magic
tech gf180mcuD
magscale 1 5
timestamp 1757618907
use signal_pad_pin  signal_pad_pin_0
timestamp 1757356153
transform 1 0 -1534 0 1 -35000
box 1534 34900 5966 35000
use signal_stub  signal_stub_0
timestamp 1757618801
transform 1 0 0 0 1 0
box 0 0 4432 800
use signal_taper  signal_taper_0
timestamp 1757356446
transform 1 0 0 0 1 800
box 0 0 4432 616
<< end >>
