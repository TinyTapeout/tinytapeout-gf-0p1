VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO loopback
  CLASS COVER ;
  FOREIGN loopback ;
  ORIGIN 0.000 0.000 ;
  SIZE 100.380 BY 0.380 ;
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 0.000 0.380 0.380 ;
    END
  END A
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 100.000 0.000 100.380 0.380 ;
    END
  END B
  OBS
      LAYER Metal2 ;
        RECT 0.380 0.000 100.000 0.380 ;
  END
END loopback
END LIBRARY

