VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_logo
  CLASS COVER ;
  FOREIGN tt_logo ;
  ORIGIN 0.000 0.000 ;
  SIZE 225.280 BY 225.280 ;
  PIN dummy
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 109.120 212.520 114.840 212.960 ;
        RECT 102.520 212.080 122.760 212.520 ;
        RECT 99.000 211.640 126.280 212.080 ;
        RECT 95.920 211.200 129.360 211.640 ;
        RECT 93.280 210.760 131.560 211.200 ;
        RECT 91.080 210.320 133.760 210.760 ;
        RECT 89.320 209.880 135.960 210.320 ;
        RECT 87.560 209.440 137.720 209.880 ;
        RECT 85.800 209.000 139.480 209.440 ;
        RECT 84.480 208.560 140.800 209.000 ;
        RECT 82.720 208.120 142.560 208.560 ;
        RECT 81.400 207.680 143.880 208.120 ;
        RECT 80.080 207.240 145.200 207.680 ;
        RECT 78.760 206.800 146.520 207.240 ;
        RECT 77.880 206.360 147.400 206.800 ;
        RECT 76.560 205.920 148.720 206.360 ;
        RECT 75.680 205.480 149.600 205.920 ;
        RECT 74.360 205.040 150.920 205.480 ;
        RECT 73.480 204.600 151.800 205.040 ;
        RECT 72.160 204.160 153.120 204.600 ;
        RECT 71.280 203.720 154.000 204.160 ;
        RECT 70.400 203.280 154.880 203.720 ;
        RECT 69.520 202.840 155.760 203.280 ;
        RECT 68.640 202.400 156.640 202.840 ;
        RECT 67.760 201.960 157.520 202.400 ;
        RECT 66.880 201.520 158.400 201.960 ;
        RECT 66.000 201.080 159.280 201.520 ;
        RECT 65.120 200.640 160.160 201.080 ;
        RECT 64.240 200.200 161.040 200.640 ;
        RECT 63.360 199.760 161.920 200.200 ;
        RECT 62.920 199.320 162.360 199.760 ;
        RECT 62.040 198.880 163.240 199.320 ;
        RECT 61.160 198.440 164.120 198.880 ;
        RECT 60.280 198.000 164.560 198.440 ;
        RECT 59.840 197.560 165.440 198.000 ;
        RECT 58.960 197.120 166.320 197.560 ;
        RECT 58.520 196.680 106.920 197.120 ;
        RECT 118.360 196.680 166.760 197.120 ;
        RECT 57.640 196.240 102.080 196.680 ;
        RECT 123.200 196.240 167.640 196.680 ;
        RECT 57.200 195.800 99.000 196.240 ;
        RECT 126.280 195.800 168.080 196.240 ;
        RECT 56.320 195.360 96.800 195.800 ;
        RECT 128.480 195.360 168.960 195.800 ;
        RECT 55.880 194.920 94.600 195.360 ;
        RECT 130.680 194.920 169.400 195.360 ;
        RECT 55.000 194.480 92.840 194.920 ;
        RECT 132.440 194.480 170.280 194.920 ;
        RECT 54.560 194.040 91.080 194.480 ;
        RECT 134.200 194.040 170.720 194.480 ;
        RECT 53.680 193.600 89.320 194.040 ;
        RECT 135.960 193.600 171.160 194.040 ;
        RECT 53.240 193.160 88.000 193.600 ;
        RECT 137.280 193.160 172.040 193.600 ;
        RECT 52.800 192.720 86.680 193.160 ;
        RECT 138.600 192.720 172.480 193.160 ;
        RECT 51.920 192.280 85.360 192.720 ;
        RECT 139.920 192.280 173.360 192.720 ;
        RECT 51.480 191.840 84.040 192.280 ;
        RECT 141.240 191.840 173.800 192.280 ;
        RECT 51.040 191.400 82.720 191.840 ;
        RECT 142.560 191.400 174.240 191.840 ;
        RECT 50.600 190.960 81.840 191.400 ;
        RECT 143.440 190.960 174.680 191.400 ;
        RECT 49.720 190.520 80.520 190.960 ;
        RECT 144.760 190.520 175.560 190.960 ;
        RECT 49.280 190.080 79.640 190.520 ;
        RECT 145.640 190.080 176.000 190.520 ;
        RECT 48.840 189.640 78.320 190.080 ;
        RECT 146.520 189.640 176.440 190.080 ;
        RECT 48.400 189.200 77.440 189.640 ;
        RECT 147.840 189.200 176.880 189.640 ;
        RECT 47.520 188.760 76.560 189.200 ;
        RECT 148.720 188.760 177.320 189.200 ;
        RECT 47.080 188.320 75.680 188.760 ;
        RECT 149.600 188.320 178.200 188.760 ;
        RECT 46.640 187.880 74.800 188.320 ;
        RECT 150.480 187.880 178.640 188.320 ;
        RECT 46.200 187.440 73.920 187.880 ;
        RECT 151.360 187.440 179.080 187.880 ;
        RECT 45.760 187.000 73.040 187.440 ;
        RECT 152.240 187.000 179.520 187.440 ;
        RECT 45.320 186.560 72.160 187.000 ;
        RECT 153.120 186.560 179.960 187.000 ;
        RECT 44.880 186.120 71.280 186.560 ;
        RECT 153.560 186.120 180.400 186.560 ;
        RECT 44.440 185.680 70.840 186.120 ;
        RECT 154.440 185.680 180.840 186.120 ;
        RECT 44.000 185.240 69.960 185.680 ;
        RECT 155.320 185.240 181.280 185.680 ;
        RECT 43.560 184.800 69.080 185.240 ;
        RECT 156.200 184.800 181.720 185.240 ;
        RECT 42.680 184.360 68.640 184.800 ;
        RECT 156.640 184.360 182.160 184.800 ;
        RECT 42.240 183.920 67.760 184.360 ;
        RECT 157.520 183.920 182.600 184.360 ;
        RECT 41.800 183.480 67.320 183.920 ;
        RECT 157.960 183.480 183.480 183.920 ;
        RECT 41.360 183.040 66.440 183.480 ;
        RECT 158.840 183.040 183.920 183.480 ;
        RECT 40.920 182.600 66.000 183.040 ;
        RECT 159.720 182.600 183.920 183.040 ;
        RECT 40.480 182.160 65.120 182.600 ;
        RECT 160.160 182.160 184.360 182.600 ;
        RECT 40.480 181.720 64.680 182.160 ;
        RECT 160.600 181.720 184.800 182.160 ;
        RECT 40.040 181.280 63.800 181.720 ;
        RECT 161.480 181.280 185.240 181.720 ;
        RECT 39.600 180.840 63.360 181.280 ;
        RECT 161.920 180.840 185.680 181.280 ;
        RECT 39.160 180.400 62.480 180.840 ;
        RECT 162.800 180.400 186.120 180.840 ;
        RECT 38.720 179.960 62.040 180.400 ;
        RECT 163.240 179.960 186.560 180.400 ;
        RECT 38.280 179.520 61.600 179.960 ;
        RECT 163.680 179.520 187.000 179.960 ;
        RECT 37.840 179.080 60.720 179.520 ;
        RECT 164.560 179.080 187.440 179.520 ;
        RECT 37.400 178.640 60.280 179.080 ;
        RECT 165.000 178.640 187.880 179.080 ;
        RECT 36.960 178.200 59.840 178.640 ;
        RECT 165.440 178.200 188.320 178.640 ;
        RECT 36.520 177.760 59.400 178.200 ;
        RECT 165.880 177.760 188.760 178.200 ;
        RECT 36.080 177.320 58.520 177.760 ;
        RECT 166.760 177.320 188.760 177.760 ;
        RECT 36.080 176.880 58.080 177.320 ;
        RECT 167.200 176.880 189.200 177.320 ;
        RECT 35.640 176.440 57.640 176.880 ;
        RECT 167.640 176.440 189.640 176.880 ;
        RECT 35.200 176.000 57.200 176.440 ;
        RECT 168.080 176.000 190.080 176.440 ;
        RECT 34.760 175.560 56.760 176.000 ;
        RECT 168.520 175.560 190.520 176.000 ;
        RECT 34.320 175.120 56.320 175.560 ;
        RECT 168.960 175.120 190.960 175.560 ;
        RECT 34.320 174.680 55.880 175.120 ;
        RECT 169.400 174.680 190.960 175.120 ;
        RECT 33.880 174.240 55.440 174.680 ;
        RECT 169.840 174.240 191.400 174.680 ;
        RECT 33.440 173.800 54.560 174.240 ;
        RECT 170.720 173.800 191.840 174.240 ;
        RECT 33.000 173.360 54.120 173.800 ;
        RECT 171.160 173.360 192.280 173.800 ;
        RECT 32.560 172.920 53.680 173.360 ;
        RECT 171.600 172.920 192.720 173.360 ;
        RECT 32.560 172.480 53.240 172.920 ;
        RECT 172.040 172.480 192.720 172.920 ;
        RECT 32.120 172.040 52.800 172.480 ;
        RECT 172.480 172.040 193.160 172.480 ;
        RECT 31.680 171.600 52.360 172.040 ;
        RECT 172.920 171.600 193.600 172.040 ;
        RECT 31.240 171.160 52.360 171.600 ;
        RECT 173.360 171.160 193.600 171.600 ;
        RECT 31.240 170.720 131.560 171.160 ;
        RECT 173.800 170.720 194.040 171.160 ;
        RECT 30.800 170.280 131.560 170.720 ;
        RECT 30.360 169.400 131.560 170.280 ;
        RECT 174.240 170.280 194.480 170.720 ;
        RECT 174.240 169.840 194.920 170.280 ;
        RECT 174.680 169.400 194.920 169.840 ;
        RECT 29.920 168.960 131.560 169.400 ;
        RECT 175.120 168.960 195.360 169.400 ;
        RECT 29.480 168.080 131.560 168.960 ;
        RECT 175.560 168.520 195.800 168.960 ;
        RECT 176.000 168.080 195.800 168.520 ;
        RECT 29.040 167.640 131.560 168.080 ;
        RECT 176.440 167.640 196.240 168.080 ;
        RECT 28.600 166.760 131.560 167.640 ;
        RECT 176.880 167.200 196.680 167.640 ;
        RECT 177.320 166.760 196.680 167.200 ;
        RECT 28.160 166.320 131.560 166.760 ;
        RECT 27.720 165.440 131.560 166.320 ;
        RECT 177.760 166.320 197.120 166.760 ;
        RECT 177.760 165.880 197.560 166.320 ;
        RECT 178.200 165.440 197.560 165.880 ;
        RECT 27.280 165.000 131.560 165.440 ;
        RECT 178.640 165.000 198.000 165.440 ;
        RECT 26.840 164.120 131.560 165.000 ;
        RECT 179.080 164.560 198.440 165.000 ;
        RECT 26.400 163.240 131.560 164.120 ;
        RECT 179.520 164.120 198.440 164.560 ;
        RECT 179.520 163.680 198.880 164.120 ;
        RECT 179.960 163.240 198.880 163.680 ;
        RECT 25.960 162.360 131.560 163.240 ;
        RECT 180.400 162.800 199.320 163.240 ;
        RECT 25.520 161.920 131.560 162.360 ;
        RECT 180.840 162.360 199.320 162.800 ;
        RECT 180.840 161.920 199.760 162.360 ;
        RECT 25.080 161.040 131.560 161.920 ;
        RECT 181.280 161.480 200.200 161.920 ;
        RECT 24.640 160.160 131.560 161.040 ;
        RECT 181.720 161.040 200.200 161.480 ;
        RECT 181.720 160.600 200.640 161.040 ;
        RECT 182.160 160.160 200.640 160.600 ;
        RECT 24.200 159.280 131.560 160.160 ;
        RECT 182.600 159.720 201.080 160.160 ;
        RECT 23.760 158.400 131.560 159.280 ;
        RECT 183.040 159.280 201.080 159.720 ;
        RECT 183.040 158.840 201.520 159.280 ;
        RECT 23.320 157.520 131.560 158.400 ;
        RECT 183.480 158.400 201.520 158.840 ;
        RECT 183.480 157.960 201.960 158.400 ;
        RECT 183.920 157.520 201.960 157.960 ;
        RECT 22.880 156.640 131.560 157.520 ;
        RECT 184.360 156.640 202.400 157.520 ;
        RECT 22.440 155.760 131.560 156.640 ;
        RECT 184.800 156.200 202.840 156.640 ;
        RECT 22.000 154.880 131.560 155.760 ;
        RECT 185.240 155.760 202.840 156.200 ;
        RECT 185.240 155.320 203.280 155.760 ;
        RECT 21.560 154.000 131.560 154.880 ;
        RECT 185.680 154.880 203.280 155.320 ;
        RECT 185.680 154.440 203.720 154.880 ;
        RECT 21.120 153.120 131.560 154.000 ;
        RECT 186.120 154.000 203.720 154.440 ;
        RECT 186.120 153.560 204.160 154.000 ;
        RECT 186.560 153.120 204.160 153.560 ;
        RECT 20.680 151.800 131.560 153.120 ;
        RECT 187.000 152.240 204.600 153.120 ;
        RECT 20.240 150.920 131.560 151.800 ;
        RECT 187.440 151.360 205.040 152.240 ;
        RECT 19.800 150.040 131.560 150.920 ;
        RECT 187.880 150.920 205.040 151.360 ;
        RECT 187.880 150.480 205.480 150.920 ;
        RECT 19.360 148.720 131.560 150.040 ;
        RECT 188.320 150.040 205.480 150.480 ;
        RECT 188.320 149.600 205.920 150.040 ;
        RECT 188.760 148.720 205.920 149.600 ;
        RECT 18.920 147.400 131.560 148.720 ;
        RECT 189.200 147.840 206.360 148.720 ;
        RECT 18.480 146.520 131.560 147.400 ;
        RECT 189.640 146.520 206.800 147.840 ;
        RECT 18.040 145.200 131.560 146.520 ;
        RECT 190.080 145.640 207.240 146.520 ;
        RECT 17.600 143.880 131.560 145.200 ;
        RECT 190.520 145.200 207.240 145.640 ;
        RECT 190.520 144.760 207.680 145.200 ;
        RECT 17.160 143.440 131.560 143.880 ;
        RECT 190.960 143.880 207.680 144.760 ;
        RECT 190.960 143.440 208.120 143.880 ;
        RECT 14.960 134.640 31.240 135.080 ;
        RECT 14.960 134.200 30.800 134.640 ;
        RECT 14.520 132.880 30.800 134.200 ;
        RECT 14.520 132.440 30.360 132.880 ;
        RECT 14.080 131.120 30.360 132.440 ;
        RECT 14.080 129.800 29.920 131.120 ;
        RECT 13.640 128.920 29.920 129.800 ;
        RECT 13.640 127.160 29.480 128.920 ;
        RECT 13.200 126.720 29.480 127.160 ;
        RECT 13.200 123.640 29.040 126.720 ;
        RECT 12.760 119.680 28.600 123.640 ;
        RECT 72.600 121.880 102.520 143.440 ;
        RECT 191.400 142.560 208.120 143.440 ;
        RECT 191.840 141.240 208.560 142.560 ;
        RECT 192.280 140.800 208.560 141.240 ;
        RECT 192.280 139.920 209.000 140.800 ;
        RECT 192.720 139.480 209.000 139.920 ;
        RECT 192.720 138.600 209.440 139.480 ;
        RECT 193.160 137.720 209.440 138.600 ;
        RECT 193.160 137.280 209.880 137.720 ;
        RECT 193.600 135.960 209.880 137.280 ;
        RECT 194.040 134.200 210.320 135.960 ;
        RECT 194.480 132.440 210.760 134.200 ;
        RECT 194.920 132.000 210.760 132.440 ;
        RECT 194.920 130.680 211.200 132.000 ;
        RECT 195.360 129.800 211.200 130.680 ;
        RECT 195.360 128.480 211.640 129.800 ;
        RECT 195.800 126.720 211.640 128.480 ;
        RECT 195.800 126.280 212.080 126.720 ;
        RECT 196.240 123.200 212.080 126.280 ;
        RECT 196.240 122.760 212.520 123.200 ;
        RECT 12.760 118.360 28.160 119.680 ;
        RECT 12.320 107.360 28.160 118.360 ;
        RECT 12.760 106.040 28.160 107.360 ;
        RECT 12.760 101.640 28.600 106.040 ;
        RECT 13.200 98.560 29.040 101.640 ;
        RECT 13.200 98.120 29.480 98.560 ;
        RECT 13.640 96.360 29.480 98.120 ;
        RECT 13.640 95.480 29.920 96.360 ;
        RECT 14.080 94.160 29.920 95.480 ;
        RECT 72.600 94.160 178.200 121.880 ;
        RECT 196.680 118.360 212.520 122.760 ;
        RECT 197.120 117.920 212.520 118.360 ;
        RECT 197.120 107.360 212.960 117.920 ;
        RECT 197.120 106.480 212.520 107.360 ;
        RECT 196.680 102.080 212.520 106.480 ;
        RECT 196.240 101.640 212.520 102.080 ;
        RECT 196.240 99.000 212.080 101.640 ;
        RECT 195.800 98.120 212.080 99.000 ;
        RECT 195.800 96.800 211.640 98.120 ;
        RECT 195.360 95.480 211.640 96.800 ;
        RECT 195.360 94.600 211.200 95.480 ;
        RECT 14.080 93.280 30.360 94.160 ;
        RECT 14.520 92.400 30.360 93.280 ;
        RECT 14.520 91.080 30.800 92.400 ;
        RECT 14.960 90.640 30.800 91.080 ;
        RECT 14.960 89.320 31.240 90.640 ;
        RECT 15.400 87.560 31.680 89.320 ;
        RECT 15.400 87.120 32.120 87.560 ;
        RECT 15.840 86.240 32.120 87.120 ;
        RECT 15.840 85.800 32.560 86.240 ;
        RECT 16.280 84.920 32.560 85.800 ;
        RECT 16.280 84.040 33.000 84.920 ;
        RECT 16.720 83.600 33.000 84.040 ;
        RECT 16.720 82.720 33.440 83.600 ;
        RECT 17.160 81.400 33.880 82.720 ;
        RECT 17.600 80.520 34.320 81.400 ;
        RECT 17.600 80.080 34.760 80.520 ;
        RECT 18.040 79.200 34.760 80.080 ;
        RECT 18.040 78.760 35.200 79.200 ;
        RECT 18.480 78.320 35.200 78.760 ;
        RECT 18.480 77.440 35.640 78.320 ;
        RECT 18.920 76.560 36.080 77.440 ;
        RECT 19.360 75.680 36.520 76.560 ;
        RECT 72.600 75.680 102.520 94.160 ;
        RECT 19.360 75.240 36.960 75.680 ;
        RECT 19.800 74.800 36.960 75.240 ;
        RECT 19.800 74.360 37.400 74.800 ;
        RECT 20.240 73.920 37.400 74.360 ;
        RECT 20.240 73.040 37.840 73.920 ;
        RECT 20.680 72.160 38.280 73.040 ;
        RECT 21.120 71.280 38.720 72.160 ;
        RECT 21.560 70.840 39.160 71.280 ;
        RECT 21.560 70.400 39.600 70.840 ;
        RECT 22.000 69.960 39.600 70.400 ;
        RECT 22.000 69.080 40.040 69.960 ;
        RECT 22.440 68.200 40.480 69.080 ;
        RECT 22.880 67.760 40.920 68.200 ;
        RECT 23.320 66.880 41.360 67.760 ;
        RECT 23.760 66.440 41.800 66.880 ;
        RECT 23.760 66.000 42.240 66.440 ;
        RECT 24.200 65.560 42.240 66.000 ;
        RECT 24.200 65.120 42.680 65.560 ;
        RECT 24.640 64.240 43.120 65.120 ;
        RECT 25.080 63.800 43.560 64.240 ;
        RECT 25.080 63.360 44.000 63.800 ;
        RECT 25.520 62.480 44.440 63.360 ;
        RECT 25.960 62.040 44.880 62.480 ;
        RECT 26.400 61.600 45.320 62.040 ;
        RECT 26.400 61.160 45.760 61.600 ;
        RECT 26.840 60.720 45.760 61.160 ;
        RECT 26.840 60.280 46.200 60.720 ;
        RECT 27.280 59.840 46.640 60.280 ;
        RECT 27.720 58.960 47.080 59.840 ;
        RECT 28.160 58.520 47.520 58.960 ;
        RECT 28.600 58.080 47.960 58.520 ;
        RECT 28.600 57.640 48.400 58.080 ;
        RECT 29.040 57.200 48.840 57.640 ;
        RECT 29.040 56.760 49.280 57.200 ;
        RECT 29.480 56.320 49.720 56.760 ;
        RECT 29.920 55.880 50.160 56.320 ;
        RECT 30.360 55.440 50.160 55.880 ;
        RECT 30.360 55.000 50.600 55.440 ;
        RECT 30.800 54.560 51.040 55.000 ;
        RECT 31.240 54.120 51.480 54.560 ;
        RECT 31.240 53.680 51.920 54.120 ;
        RECT 31.680 53.240 52.360 53.680 ;
        RECT 32.120 52.800 52.800 53.240 ;
        RECT 32.560 52.360 53.240 52.800 ;
        RECT 32.560 51.920 53.680 52.360 ;
        RECT 33.000 51.480 54.120 51.920 ;
        RECT 33.440 51.040 54.560 51.480 ;
        RECT 33.880 50.600 55.000 51.040 ;
        RECT 33.880 50.160 55.440 50.600 ;
        RECT 34.320 49.720 56.320 50.160 ;
        RECT 34.760 49.280 56.760 49.720 ;
        RECT 35.200 48.840 57.200 49.280 ;
        RECT 35.640 48.400 57.640 48.840 ;
        RECT 36.080 47.960 58.080 48.400 ;
        RECT 36.080 47.520 58.520 47.960 ;
        RECT 36.520 47.080 59.400 47.520 ;
        RECT 36.960 46.640 59.840 47.080 ;
        RECT 37.400 46.200 60.280 46.640 ;
        RECT 37.840 45.760 60.720 46.200 ;
        RECT 38.280 45.320 61.600 45.760 ;
        RECT 38.720 44.880 62.040 45.320 ;
        RECT 39.160 44.440 62.480 44.880 ;
        RECT 39.600 44.000 63.360 44.440 ;
        RECT 39.600 43.560 63.800 44.000 ;
        RECT 40.040 43.120 64.240 43.560 ;
        RECT 40.480 42.680 65.120 43.120 ;
        RECT 40.920 42.240 65.560 42.680 ;
        RECT 41.360 41.800 66.440 42.240 ;
        RECT 41.800 41.360 66.880 41.800 ;
        RECT 42.240 40.920 67.760 41.360 ;
        RECT 42.680 40.480 68.640 40.920 ;
        RECT 43.120 40.040 69.080 40.480 ;
        RECT 44.000 39.600 69.960 40.040 ;
        RECT 44.440 39.160 70.840 39.600 ;
        RECT 44.880 38.720 71.280 39.160 ;
        RECT 45.320 38.280 72.160 38.720 ;
        RECT 45.760 37.840 73.040 38.280 ;
        RECT 46.200 37.400 73.920 37.840 ;
        RECT 46.640 36.960 74.800 37.400 ;
        RECT 47.080 36.520 75.680 36.960 ;
        RECT 47.520 36.080 76.560 36.520 ;
        RECT 48.400 35.640 77.440 36.080 ;
        RECT 48.840 35.200 78.320 35.640 ;
        RECT 49.280 34.760 79.640 35.200 ;
        RECT 49.720 34.320 80.520 34.760 ;
        RECT 50.600 33.880 81.840 34.320 ;
        RECT 51.040 33.440 82.720 33.880 ;
        RECT 51.480 33.000 84.040 33.440 ;
        RECT 51.920 32.560 85.360 33.000 ;
        RECT 52.800 32.120 86.680 32.560 ;
        RECT 53.240 31.680 88.000 32.120 ;
        RECT 53.680 31.240 89.320 31.680 ;
        RECT 54.560 30.800 91.080 31.240 ;
        RECT 55.000 30.360 92.840 30.800 ;
        RECT 55.880 29.920 94.600 30.360 ;
        RECT 56.320 29.480 96.800 29.920 ;
        RECT 57.200 29.040 99.000 29.480 ;
        RECT 57.640 28.600 102.080 29.040 ;
        RECT 119.240 28.600 149.160 94.160 ;
        RECT 194.920 93.280 211.200 94.600 ;
        RECT 194.920 92.840 210.760 93.280 ;
        RECT 194.480 91.080 210.760 92.840 ;
        RECT 194.040 89.320 210.320 91.080 ;
        RECT 193.600 88.880 210.320 89.320 ;
        RECT 193.600 88.000 209.880 88.880 ;
        RECT 193.160 87.120 209.880 88.000 ;
        RECT 193.160 86.680 209.440 87.120 ;
        RECT 192.720 85.800 209.440 86.680 ;
        RECT 192.720 85.360 209.000 85.800 ;
        RECT 192.280 84.040 209.000 85.360 ;
        RECT 191.840 82.720 208.560 84.040 ;
        RECT 191.400 81.840 208.120 82.720 ;
        RECT 190.960 81.400 208.120 81.840 ;
        RECT 190.960 80.520 207.680 81.400 ;
        RECT 190.520 80.080 207.680 80.520 ;
        RECT 190.520 79.640 207.240 80.080 ;
        RECT 190.080 78.760 207.240 79.640 ;
        RECT 190.080 78.320 206.800 78.760 ;
        RECT 189.640 77.440 206.800 78.320 ;
        RECT 189.200 76.560 206.360 77.440 ;
        RECT 188.760 75.680 205.920 76.560 ;
        RECT 188.320 75.240 205.920 75.680 ;
        RECT 188.320 74.800 205.480 75.240 ;
        RECT 187.880 74.360 205.480 74.800 ;
        RECT 187.880 73.920 205.040 74.360 ;
        RECT 187.440 73.040 205.040 73.920 ;
        RECT 187.000 72.160 204.600 73.040 ;
        RECT 186.560 71.280 204.160 72.160 ;
        RECT 186.120 70.840 203.720 71.280 ;
        RECT 185.680 70.400 203.720 70.840 ;
        RECT 185.680 69.960 203.280 70.400 ;
        RECT 185.240 69.080 203.280 69.960 ;
        RECT 184.800 68.640 202.840 69.080 ;
        RECT 184.360 68.200 202.840 68.640 ;
        RECT 184.360 67.760 202.400 68.200 ;
        RECT 183.920 67.320 202.400 67.760 ;
        RECT 183.920 66.880 201.960 67.320 ;
        RECT 183.480 66.440 201.960 66.880 ;
        RECT 183.040 65.560 201.520 66.440 ;
        RECT 182.600 65.120 201.080 65.560 ;
        RECT 182.160 64.680 200.640 65.120 ;
        RECT 181.720 64.240 200.640 64.680 ;
        RECT 181.720 63.800 200.200 64.240 ;
        RECT 181.280 63.360 200.200 63.800 ;
        RECT 180.840 62.480 199.760 63.360 ;
        RECT 180.400 62.040 199.320 62.480 ;
        RECT 179.960 61.600 198.880 62.040 ;
        RECT 179.520 61.160 198.880 61.600 ;
        RECT 179.520 60.720 198.440 61.160 ;
        RECT 179.080 60.280 198.440 60.720 ;
        RECT 178.640 59.840 198.000 60.280 ;
        RECT 178.200 59.400 197.560 59.840 ;
        RECT 177.760 58.960 197.560 59.400 ;
        RECT 177.760 58.520 197.120 58.960 ;
        RECT 177.320 58.080 197.120 58.520 ;
        RECT 176.880 57.640 196.680 58.080 ;
        RECT 176.440 57.200 196.240 57.640 ;
        RECT 176.000 56.760 196.240 57.200 ;
        RECT 175.560 56.320 195.800 56.760 ;
        RECT 175.120 55.880 195.360 56.320 ;
        RECT 174.680 55.440 195.360 55.880 ;
        RECT 174.680 55.000 194.920 55.440 ;
        RECT 174.240 54.560 194.480 55.000 ;
        RECT 173.800 54.120 194.040 54.560 ;
        RECT 173.360 53.680 194.040 54.120 ;
        RECT 172.920 53.240 193.600 53.680 ;
        RECT 172.480 52.800 193.160 53.240 ;
        RECT 172.040 52.360 192.720 52.800 ;
        RECT 171.600 51.920 192.720 52.360 ;
        RECT 171.160 51.480 192.280 51.920 ;
        RECT 170.720 51.040 191.840 51.480 ;
        RECT 170.280 50.600 191.400 51.040 ;
        RECT 169.400 50.160 191.400 50.600 ;
        RECT 168.960 49.720 190.960 50.160 ;
        RECT 168.520 49.280 190.520 49.720 ;
        RECT 168.080 48.840 190.080 49.280 ;
        RECT 167.640 48.400 189.640 48.840 ;
        RECT 167.200 47.960 189.640 48.400 ;
        RECT 166.760 47.520 189.200 47.960 ;
        RECT 165.880 47.080 188.760 47.520 ;
        RECT 165.440 46.640 188.320 47.080 ;
        RECT 165.000 46.200 187.880 46.640 ;
        RECT 164.560 45.760 187.440 46.200 ;
        RECT 163.680 45.320 187.000 45.760 ;
        RECT 163.240 44.880 186.560 45.320 ;
        RECT 162.800 44.440 186.120 44.880 ;
        RECT 161.920 44.000 186.120 44.440 ;
        RECT 161.480 43.560 185.680 44.000 ;
        RECT 161.040 43.120 185.240 43.560 ;
        RECT 160.160 42.680 184.800 43.120 ;
        RECT 159.720 42.240 184.360 42.680 ;
        RECT 158.840 41.800 183.920 42.240 ;
        RECT 158.400 41.360 183.480 41.800 ;
        RECT 58.520 28.160 106.920 28.600 ;
        RECT 118.360 28.160 149.160 28.600 ;
        RECT 58.960 27.720 149.160 28.160 ;
        RECT 59.840 27.280 149.160 27.720 ;
        RECT 60.280 26.840 149.160 27.280 ;
        RECT 61.160 26.400 149.160 26.840 ;
        RECT 62.040 25.960 149.160 26.400 ;
        RECT 62.920 25.520 149.160 25.960 ;
        RECT 63.360 25.080 149.160 25.520 ;
        RECT 64.240 24.640 149.160 25.080 ;
        RECT 65.120 24.200 149.160 24.640 ;
        RECT 66.000 23.760 149.160 24.200 ;
        RECT 66.880 23.320 149.160 23.760 ;
        RECT 157.520 40.920 183.040 41.360 ;
        RECT 157.520 40.480 182.600 40.920 ;
        RECT 157.520 40.040 182.160 40.480 ;
        RECT 157.520 39.600 181.720 40.040 ;
        RECT 157.520 39.160 181.280 39.600 ;
        RECT 157.520 38.720 180.840 39.160 ;
        RECT 157.520 38.280 179.960 38.720 ;
        RECT 157.520 37.840 179.520 38.280 ;
        RECT 157.520 37.400 179.080 37.840 ;
        RECT 157.520 36.960 178.640 37.400 ;
        RECT 157.520 36.520 178.200 36.960 ;
        RECT 157.520 36.080 177.760 36.520 ;
        RECT 157.520 35.640 177.320 36.080 ;
        RECT 157.520 35.200 176.440 35.640 ;
        RECT 157.520 34.760 176.000 35.200 ;
        RECT 157.520 34.320 175.560 34.760 ;
        RECT 157.520 33.880 175.120 34.320 ;
        RECT 157.520 33.440 174.240 33.880 ;
        RECT 157.520 33.000 173.800 33.440 ;
        RECT 157.520 32.560 173.360 33.000 ;
        RECT 157.520 32.120 172.480 32.560 ;
        RECT 157.520 31.680 172.040 32.120 ;
        RECT 157.520 31.240 171.600 31.680 ;
        RECT 157.520 30.800 170.720 31.240 ;
        RECT 157.520 30.360 170.280 30.800 ;
        RECT 157.520 29.920 169.840 30.360 ;
        RECT 157.520 29.480 168.960 29.920 ;
        RECT 157.520 29.040 168.520 29.480 ;
        RECT 157.520 28.600 167.640 29.040 ;
        RECT 157.520 28.160 167.200 28.600 ;
        RECT 157.520 27.720 166.320 28.160 ;
        RECT 157.520 27.280 165.440 27.720 ;
        RECT 157.520 26.840 165.000 27.280 ;
        RECT 157.520 26.400 164.120 26.840 ;
        RECT 157.520 25.960 163.240 26.400 ;
        RECT 157.520 25.520 162.800 25.960 ;
        RECT 157.520 25.080 161.920 25.520 ;
        RECT 157.520 24.640 161.040 25.080 ;
        RECT 157.520 24.200 160.160 24.640 ;
        RECT 157.520 23.760 159.280 24.200 ;
        RECT 157.520 23.320 158.840 23.760 ;
        RECT 67.760 22.880 149.160 23.320 ;
        RECT 68.640 22.440 149.160 22.880 ;
        RECT 69.520 22.000 149.160 22.440 ;
        RECT 70.400 21.560 149.160 22.000 ;
        RECT 71.280 21.120 149.160 21.560 ;
        RECT 72.160 20.680 149.160 21.120 ;
        RECT 73.040 20.240 149.160 20.680 ;
        RECT 74.360 19.800 149.160 20.240 ;
        RECT 75.240 19.360 149.160 19.800 ;
        RECT 76.560 18.920 148.720 19.360 ;
        RECT 77.880 18.480 147.400 18.920 ;
        RECT 78.760 18.040 146.520 18.480 ;
        RECT 80.080 17.600 145.200 18.040 ;
        RECT 81.400 17.160 143.880 17.600 ;
        RECT 82.720 16.720 142.560 17.160 ;
        RECT 84.480 16.280 140.800 16.720 ;
        RECT 85.800 15.840 139.480 16.280 ;
        RECT 87.560 15.400 137.720 15.840 ;
        RECT 89.320 14.960 135.960 15.400 ;
        RECT 91.080 14.520 133.760 14.960 ;
        RECT 93.280 14.080 131.560 14.520 ;
        RECT 95.920 13.640 129.360 14.080 ;
        RECT 99.000 13.200 126.280 13.640 ;
        RECT 102.520 12.760 122.760 13.200 ;
        RECT 109.120 12.320 116.160 12.760 ;
    END
  END dummy
END tt_logo
END LIBRARY

