magic
tech gf180mcuD
magscale 1 10
timestamp 1757360064
<< metal2 >>
rect 127400 518884 127720 520164
rect 127400 518564 144720 518884
rect 144400 509872 144720 518564
rect 147400 510532 147720 520164
rect 147390 510212 147400 510532
rect 147720 510212 147730 510532
rect 144390 509552 144400 509872
rect 144720 509552 144730 509872
rect 74956 467400 76556 467720
rect 76236 450720 76556 467400
rect 187060 454984 188060 520444
rect 207522 518260 207598 519940
rect 227522 518660 227598 519940
rect 247522 519060 247598 519940
rect 267522 519460 267598 519940
rect 282337 519460 282413 521060
rect 267522 519384 282413 519460
rect 293940 519060 294016 521060
rect 247522 518984 294016 519060
rect 294086 518660 294162 521060
rect 227522 518584 294162 518660
rect 294232 518260 294308 521060
rect 407060 518544 408060 520444
rect 207522 518184 294308 518260
rect 405673 517544 408060 518544
rect 187050 453984 187060 454984
rect 188060 453984 188070 454984
rect 405673 453584 406673 517544
rect 427060 515544 428060 520444
rect 467400 518884 467720 520164
rect 408673 514544 428060 515544
rect 450400 518564 467720 518884
rect 408673 454984 409673 514544
rect 450400 510532 450720 518564
rect 450390 510212 450400 510532
rect 450720 510212 450730 510532
rect 518564 467400 520164 467720
rect 408663 453984 408673 454984
rect 409673 453984 409683 454984
rect 405663 452584 405673 453584
rect 406673 452584 406683 453584
rect 84244 450720 84564 450730
rect 76236 450400 84244 450720
rect 84244 450390 84564 450400
rect 510000 450720 510320 450730
rect 518564 450720 518884 467400
rect 510320 450400 518884 450720
rect 510000 450390 510320 450400
rect 510660 447720 510980 447730
rect 510980 447400 520164 447720
rect 510660 447390 510980 447400
rect 74676 427060 80576 428060
rect 79576 409673 80576 427060
rect 139640 409673 140640 409683
rect 79576 408673 139640 409673
rect 139640 408663 140640 408673
rect 454544 408060 455544 408070
rect 74676 407060 77576 408060
rect 76576 406673 77576 407060
rect 455544 407060 520444 408060
rect 454544 407050 455544 407060
rect 141040 406673 142040 406683
rect 76576 405673 141040 406673
rect 141040 405663 142040 405673
rect 453144 189447 454144 189457
rect 454144 188447 518544 189447
rect 453144 188437 454144 188447
rect 139640 188060 140640 188070
rect 74676 187060 139640 188060
rect 517544 188060 518544 188447
rect 517544 187060 520444 188060
rect 139640 187050 140640 187060
rect 454544 186447 455544 186457
rect 455544 185447 515544 186447
rect 454544 185437 455544 185447
rect 514544 168060 515544 185447
rect 514544 167060 520444 168060
rect 84244 147720 84564 147730
rect 74956 147400 84244 147720
rect 84244 147390 84564 147400
rect 84904 144720 85224 144730
rect 76236 144400 84904 144720
rect 76236 127720 76556 144400
rect 84904 144390 85224 144400
rect 510660 144720 510980 144730
rect 510980 144400 518884 144720
rect 510660 144390 510980 144400
rect 188437 141488 188447 142488
rect 189447 141488 189457 142488
rect 185437 140088 185447 141088
rect 186447 140088 186457 141088
rect 74956 127400 76556 127720
rect 144390 84244 144400 84564
rect 144720 84244 144730 84564
rect 144400 76556 144720 84244
rect 185447 80576 186447 140088
rect 127400 76236 144720 76556
rect 167060 79576 186447 80576
rect 127400 74956 127720 76236
rect 167060 74676 168060 79576
rect 188447 77576 189447 141488
rect 407050 140088 407060 141088
rect 408060 140088 408070 141088
rect 187060 76576 189447 77576
rect 187060 74676 188060 76576
rect 207522 75180 207598 76136
rect 227522 75180 227598 76136
rect 407060 74676 408060 140088
rect 518564 127720 518884 144400
rect 518564 127400 520164 127720
rect 450390 85690 450400 86010
rect 450720 85690 450730 86010
rect 447390 85030 447400 85350
rect 447720 85030 447730 85350
rect 447400 74956 447720 85030
rect 450400 76556 450720 85690
rect 450400 76236 467720 76556
rect 467400 74956 467720 76236
<< via2 >>
rect 147400 510212 147720 510532
rect 144400 509552 144720 509872
rect 187060 453984 188060 454984
rect 450400 510212 450720 510532
rect 408673 453984 409673 454984
rect 405673 452584 406673 453584
rect 84244 450400 84564 450720
rect 510000 450400 510320 450720
rect 510660 447400 510980 447720
rect 139640 408673 140640 409673
rect 454544 407060 455544 408060
rect 141040 405673 142040 406673
rect 453144 188447 454144 189447
rect 139640 187060 140640 188060
rect 454544 185447 455544 186447
rect 84244 147400 84564 147720
rect 84904 144400 85224 144720
rect 510660 144400 510980 144720
rect 188447 141488 189447 142488
rect 185447 140088 186447 141088
rect 144400 84244 144720 84564
rect 407060 140088 408060 141088
rect 450400 85690 450720 86010
rect 447400 85030 447720 85350
<< metal3 >>
rect 147400 510532 147720 510541
rect 450400 510532 450720 510541
rect 147391 510212 147400 510532
rect 147720 510212 147729 510532
rect 450391 510212 450400 510532
rect 450720 510212 450729 510532
rect 147400 510203 147720 510212
rect 450400 510203 450720 510212
rect 144400 509872 144720 509881
rect 144391 509552 144400 509872
rect 144720 509552 144729 509872
rect 144400 509543 144720 509552
rect 187060 454984 188060 454993
rect 408673 454984 409673 454993
rect 187051 453984 187060 454984
rect 188060 453984 188069 454984
rect 408664 453984 408673 454984
rect 409673 453984 409682 454984
rect 187060 453975 188060 453984
rect 408673 453975 409673 453984
rect 405673 453584 406673 453593
rect 405664 452584 405673 453584
rect 406673 452584 406682 453584
rect 405673 452575 406673 452584
rect 84244 450720 84564 450729
rect 510000 450720 510320 450729
rect 84235 450400 84244 450720
rect 84564 450400 84573 450720
rect 509991 450400 510000 450720
rect 510320 450400 510329 450720
rect 84244 450391 84564 450400
rect 510000 450391 510320 450400
rect 510660 447720 510980 447729
rect 510651 447400 510660 447720
rect 510980 447400 510989 447720
rect 510660 447391 510980 447400
rect 139640 409673 140640 409682
rect 139631 408673 139640 409673
rect 140640 408673 140649 409673
rect 139640 408664 140640 408673
rect 454544 408060 455544 408069
rect 454535 407060 454544 408060
rect 455544 407060 455553 408060
rect 454544 407051 455544 407060
rect 141040 406673 142040 406682
rect 141031 405673 141040 406673
rect 142040 405673 142049 406673
rect 141040 405664 142040 405673
rect 453144 189447 454144 189456
rect 453135 188447 453144 189447
rect 454144 188447 454153 189447
rect 453144 188438 454144 188447
rect 139640 188060 140640 188069
rect 139631 187060 139640 188060
rect 140640 187060 140649 188060
rect 139640 187051 140640 187060
rect 454544 186447 455544 186456
rect 454535 185447 454544 186447
rect 455544 185447 455553 186447
rect 454544 185438 455544 185447
rect 84244 147720 84564 147729
rect 84235 147400 84244 147720
rect 84564 147400 84573 147720
rect 84244 147391 84564 147400
rect 84904 144720 85224 144729
rect 510660 144720 510980 144729
rect 84895 144400 84904 144720
rect 85224 144400 85233 144720
rect 510651 144400 510660 144720
rect 510980 144400 510989 144720
rect 84904 144391 85224 144400
rect 510660 144391 510980 144400
rect 188447 142488 189447 142497
rect 188438 141488 188447 142488
rect 189447 141488 189456 142488
rect 188447 141479 189447 141488
rect 185447 141088 186447 141097
rect 407060 141088 408060 141097
rect 185438 140088 185447 141088
rect 186447 140088 186456 141088
rect 407051 140088 407060 141088
rect 408060 140088 408069 141088
rect 185447 140079 186447 140088
rect 407060 140079 408060 140088
rect 450400 86010 450720 86019
rect 450391 85690 450400 86010
rect 450720 85690 450729 86010
rect 450400 85681 450720 85690
rect 447400 85350 447720 85359
rect 447391 85030 447400 85350
rect 447720 85030 447729 85350
rect 447400 85021 447720 85030
rect 144400 84564 144720 84573
rect 144391 84244 144400 84564
rect 144720 84244 144729 84564
rect 144400 84235 144720 84244
<< via3 >>
rect 147400 510212 147720 510532
rect 450400 510212 450720 510532
rect 144400 509552 144720 509872
rect 187060 453984 188060 454984
rect 408673 453984 409673 454984
rect 405673 452584 406673 453584
rect 84244 450400 84564 450720
rect 510000 450400 510320 450720
rect 510660 447400 510980 447720
rect 139640 408673 140640 409673
rect 454544 407060 455544 408060
rect 141040 405673 142040 406673
rect 453144 188447 454144 189447
rect 139640 187060 140640 188060
rect 454544 185447 455544 186447
rect 84244 147400 84564 147720
rect 84904 144400 85224 144720
rect 510660 144400 510980 144720
rect 188447 141488 189447 142488
rect 185447 140088 186447 141088
rect 407060 140088 408060 141088
rect 450400 85690 450720 86010
rect 447400 85030 447720 85350
rect 144400 84244 144720 84564
<< metal4 >>
rect 147400 510532 147720 510541
rect 450400 510532 450720 510541
rect 147391 510212 147400 510532
rect 147720 510212 147729 510532
rect 450391 510212 450400 510532
rect 450720 510212 450729 510532
rect 147400 510203 147720 510212
rect 450400 510203 450720 510212
rect 144400 509872 144720 509881
rect 144391 509552 144400 509872
rect 144720 509552 144729 509872
rect 144400 509543 144720 509552
rect 187060 454984 188060 454993
rect 408673 454984 409673 454993
rect 187051 453984 187060 454984
rect 188060 453984 188069 454984
rect 408664 453984 408673 454984
rect 409673 453984 409682 454984
rect 187060 453975 188060 453984
rect 408673 453975 409673 453984
rect 405673 453584 406673 453593
rect 405664 452584 405673 453584
rect 406673 452584 406682 453584
rect 405673 452575 406673 452584
rect 84244 450720 84564 452000
rect 84235 450400 84244 450720
rect 84564 450400 84573 450720
rect 84244 449120 84564 450400
rect 84904 449120 85224 452000
rect 510000 450720 510320 452000
rect 509991 450400 510000 450720
rect 510320 450400 510329 450720
rect 510000 446120 510320 450400
rect 510660 447720 510980 452000
rect 510651 447400 510660 447720
rect 510980 447400 510989 447720
rect 510660 446120 510980 447400
rect 139640 409673 140640 413673
rect 139631 408673 139640 409673
rect 140640 408673 140649 409673
rect 139640 401673 140640 408673
rect 141040 406673 142040 413673
rect 141031 405673 141040 406673
rect 142040 405673 142049 406673
rect 141040 401673 142040 405673
rect 453144 403060 454144 412060
rect 454544 408060 455544 412060
rect 454535 407060 454544 408060
rect 455544 407060 455553 408060
rect 454544 403060 455544 407060
rect 139640 188060 140640 192060
rect 139631 187060 139640 188060
rect 140640 187060 140649 188060
rect 139640 183060 140640 187060
rect 141040 183060 142040 192060
rect 453144 189447 454144 193447
rect 453135 188447 453144 189447
rect 454144 188447 454153 189447
rect 453144 181447 454144 188447
rect 454544 186447 455544 193447
rect 454535 185447 454544 186447
rect 455544 185447 455553 186447
rect 454544 181447 455544 185447
rect 84244 147720 84564 149000
rect 84235 147400 84244 147720
rect 84564 147400 84573 147720
rect 84244 143120 84564 147400
rect 84904 144720 85224 149000
rect 84895 144400 84904 144720
rect 85224 144400 85233 144720
rect 84904 143120 85224 144400
rect 510000 143120 510320 146000
rect 510660 144720 510980 146000
rect 510651 144400 510660 144720
rect 510980 144400 510989 144720
rect 510660 143120 510980 144400
rect 188447 142488 189447 142497
rect 188438 141488 188447 142488
rect 189447 141488 189456 142488
rect 188447 141479 189447 141488
rect 185447 141088 186447 141097
rect 407060 141088 408060 141097
rect 185438 140088 185447 141088
rect 186447 140088 186456 141088
rect 407051 140088 407060 141088
rect 408060 140088 408069 141088
rect 185447 140079 186447 140088
rect 407060 140079 408060 140088
rect 450400 86010 450720 86019
rect 450391 85690 450400 86010
rect 450720 85690 450729 86010
rect 450400 85681 450720 85690
rect 447400 85350 447720 85359
rect 447391 85030 447400 85350
rect 447720 85030 447729 85350
rect 447400 85021 447720 85030
rect 144400 84564 144720 84573
rect 144391 84244 144400 84564
rect 144720 84244 144729 84564
rect 144400 84235 144720 84244
<< via4 >>
rect 147400 510212 147720 510532
rect 450400 510212 450720 510532
rect 144400 509552 144720 509872
rect 187060 453984 188060 454984
rect 408673 453984 409673 454984
rect 405673 452584 406673 453584
rect 188447 141488 189447 142488
rect 185447 140088 186447 141088
rect 407060 140088 408060 141088
rect 450400 85690 450720 86010
rect 447400 85030 447720 85350
rect 144400 84244 144720 84564
<< metal5 >>
rect 147400 510532 147720 510541
rect 450400 510532 450720 510541
rect 143120 510212 147400 510532
rect 147720 510212 149000 510532
rect 449120 510212 450400 510532
rect 450720 510212 452000 510532
rect 147400 510203 147720 510212
rect 450400 510203 450720 510212
rect 144400 509872 144720 509881
rect 143120 509552 144400 509872
rect 144720 509552 149000 509872
rect 449120 509552 452000 509872
rect 144400 509543 144720 509552
rect 187060 454984 188060 454993
rect 408673 454984 409673 454993
rect 183060 453984 187060 454984
rect 188060 453984 192060 454984
rect 401673 453984 408673 454984
rect 409673 453984 413673 454984
rect 187060 453975 188060 453984
rect 408673 453975 409673 453984
rect 405673 453584 406673 453593
rect 183060 452584 192060 453584
rect 401673 452584 405673 453584
rect 406673 452584 413673 453584
rect 405673 452575 406673 452584
rect 188447 142488 189447 142497
rect 181447 141488 188447 142488
rect 189447 141488 193447 142488
rect 403060 141488 412060 142488
rect 188447 141479 189447 141488
rect 185447 141088 186447 141097
rect 407060 141088 408060 141097
rect 181447 140088 185447 141088
rect 186447 140088 193447 141088
rect 403060 140088 407060 141088
rect 408060 140088 412060 141088
rect 185447 140079 186447 140088
rect 407060 140079 408060 140088
rect 450400 86010 450720 86019
rect 446120 85690 450400 86010
rect 450720 85690 452000 86010
rect 450400 85681 450720 85690
rect 447400 85350 447720 85359
rect 143120 84904 146000 85224
rect 446120 85030 447400 85350
rect 447720 85030 452000 85350
rect 447400 85021 447720 85030
rect 144400 84564 144720 84573
rect 143120 84244 144400 84564
rect 144720 84244 146000 84564
rect 144400 84235 144720 84244
use power_taper  power_taper_0
timestamp 1757356513
transform 1 0 120332 0 1 74060
box 0 -200 14456 1344
use power_taper  power_taper_2
timestamp 1757356513
transform 1 0 160332 0 1 74060
box 0 -200 14456 1344
use power_taper  power_taper_3
timestamp 1757356513
transform 1 0 180332 0 1 74060
box 0 -200 14456 1344
use power_taper  power_taper_4
timestamp 1757356513
transform 1 0 400332 0 1 74060
box 0 -200 14456 1344
use power_taper  power_taper_6
timestamp 1757356513
transform 1 0 440332 0 1 74060
box 0 -200 14456 1344
use power_taper  power_taper_7
timestamp 1757356513
transform 1 0 460332 0 1 74060
box 0 -200 14456 1344
use power_taper  power_taper_8
timestamp 1757356513
transform 0 -1 521060 1 0 120332
box 0 -200 14456 1344
use power_taper  power_taper_10
timestamp 1757356513
transform 0 -1 521060 1 0 160332
box 0 -200 14456 1344
use power_taper  power_taper_11
timestamp 1757356513
transform 0 -1 521060 1 0 180332
box 0 -200 14456 1344
use power_taper  power_taper_12
timestamp 1757356513
transform 0 -1 521060 1 0 400332
box 0 -200 14456 1344
use power_taper  power_taper_14
timestamp 1757356513
transform 0 -1 521060 1 0 440332
box 0 -200 14456 1344
use power_taper  power_taper_15
timestamp 1757356513
transform 0 -1 521060 1 0 460332
box 0 -200 14456 1344
use power_taper  power_taper_16
timestamp 1757356513
transform -1 0 474788 0 -1 521060
box 0 -200 14456 1344
use power_taper  power_taper_18
timestamp 1757356513
transform -1 0 434788 0 -1 521060
box 0 -200 14456 1344
use power_taper  power_taper_19
timestamp 1757356513
transform -1 0 414788 0 -1 521060
box 0 -200 14456 1344
use power_taper  power_taper_20
timestamp 1757356513
transform -1 0 194788 0 -1 521060
box 0 -200 14456 1344
use power_taper  power_taper_22
timestamp 1757356513
transform -1 0 154788 0 -1 521060
box 0 -200 14456 1344
use power_taper  power_taper_23
timestamp 1757356513
transform -1 0 134788 0 -1 521060
box 0 -200 14456 1344
use power_taper  power_taper_24
timestamp 1757356513
transform 0 1 74060 -1 0 474788
box 0 -200 14456 1344
use power_taper  power_taper_26
timestamp 1757356513
transform 0 1 74060 -1 0 434788
box 0 -200 14456 1344
use power_taper  power_taper_27
timestamp 1757356513
transform 0 1 74060 -1 0 414788
box 0 -200 14456 1344
use power_taper  power_taper_28
timestamp 1757356513
transform 0 1 74060 -1 0 194788
box 0 -200 14456 1344
use power_taper  power_taper_30
timestamp 1757356513
transform 0 1 74060 -1 0 154788
box 0 -200 14456 1344
use power_taper  power_taper_31
timestamp 1757356513
transform 0 1 74060 -1 0 134788
box 0 -200 14456 1344
use signal_taper  signal_taper_0
timestamp 1757356446
transform 1 0 203128 0 1 74060
box 0 -200 8864 1232
use signal_taper  signal_taper_1
timestamp 1757356446
transform 1 0 223128 0 1 74060
box 0 -200 8864 1232
use signal_taper  signal_taper_2
timestamp 1757356446
transform -1 0 271992 0 -1 521060
box 0 -200 8864 1232
use signal_taper  signal_taper_3
timestamp 1757356446
transform -1 0 251992 0 -1 521060
box 0 -200 8864 1232
use signal_taper  signal_taper_4
timestamp 1757356446
transform -1 0 231992 0 -1 521060
box 0 -200 8864 1232
use signal_taper  signal_taper_5
timestamp 1757356446
transform -1 0 211992 0 -1 521060
box 0 -200 8864 1232
<< labels >>
flabel metal5 143120 84244 146000 84564 0 FreeSans 1024 0 0 0 vss_pad_s_2
port 1 nsew ground bidirectional
flabel metal5 181447 140088 193447 141088 0 FreeSans 1024 0 0 0 vss_pad_s_4
port 2 nsew ground bidirectional
flabel metal5 181447 141488 193447 142488 0 FreeSans 1024 0 0 0 vddcore0_pad_s_5
port 3 nsew power bidirectional
flabel metal5 403060 140088 412060 141088 0 FreeSans 1024 0 0 0 vss_pad_s_16
port 4 nsew ground bidirectional
flabel metal5 446120 85030 452000 85350 0 FreeSans 1024 0 0 0 vss_pad_s_18
port 5 nsew ground bidirectional
flabel metal5 446120 85690 452000 86010 0 FreeSans 1024 0 0 0 vddcore3_pad_s_19
port 6 nsew power bidirectional
flabel metal4 510660 143120 510980 146000 0 FreeSans 1024 90 0 0 vss_pad_e_2
port 7 nsew ground bidirectional
flabel metal4 454544 181447 455544 193447 0 FreeSans 1024 90 0 0 vss_pad_e_4
port 8 nsew ground bidirectional
flabel metal4 453144 181447 454144 193447 0 FreeSans 1024 90 0 0 vddcore0_pad_e_5
port 9 nsew power bidirectional
flabel metal4 454544 403060 455544 412060 0 FreeSans 1024 90 0 0 vss_pad_e_16
port 10 nsew ground bidirectional
flabel metal4 510660 446120 510980 452000 0 FreeSans 1024 90 0 0 vss_pad_e_18
port 11 nsew ground bidirectional
flabel metal4 510000 446120 510320 452000 0 FreeSans 1024 90 0 0 vddcore4_pad_e_19
port 12 nsew power bidirectional
flabel metal5 449120 510212 452000 510532 0 FreeSans 1024 0 0 0 vss_pad_n_2
port 13 nsew ground bidirectional
flabel metal5 401673 453984 413673 454984 0 FreeSans 1024 0 0 0 vss_pad_n_4
port 14 nsew ground bidirectional
flabel metal5 401673 452584 413673 453584 0 FreeSans 1024 0 0 0 vddcore0_pad_n_5
port 15 nsew power bidirectional
flabel metal5 183060 453984 192060 454984 0 FreeSans 1024 0 0 0 vss_pad_n_16
port 16 nsew ground bidirectional
flabel metal5 143120 510212 149000 510532 0 FreeSans 1024 0 0 0 vss_pad_n_18
port 17 nsew ground bidirectional
flabel metal5 143120 509552 149000 509872 0 FreeSans 1024 0 0 0 vddcore1_pad_n_19
port 18 nsew power bidirectional
flabel metal4 84244 449120 84564 452000 0 FreeSans 1024 90 0 0 vss_pad_w_2
port 19 nsew ground bidirectional
flabel metal4 139640 401673 140640 413673 0 FreeSans 1024 90 0 0 vss_pad_w_4
port 20 nsew ground bidirectional
flabel metal4 141040 401673 142040 413673 0 FreeSans 1024 90 0 0 vddcore0_pad_w_5
port 21 nsew power bidirectional
flabel metal4 139640 183060 140640 192060 0 FreeSans 1024 90 0 0 vss_pad_w_16
port 22 nsew ground bidirectional
flabel metal4 84244 143120 84564 149000 0 FreeSans 1024 90 0 0 vss_pad_w_18
port 23 nsew ground bidirectional
flabel metal4 84904 143120 85224 149000 0 FreeSans 1024 90 0 0 vddcore2_pad_w_19
port 24 nsew power bidirectional
flabel metal2 207522 75180 207598 76136 0 FreeSans 1024 0 0 0 loop_pad_s_6
port 25 nsew signal bidirectional
flabel metal2 227522 75180 227598 76136 0 FreeSans 1024 0 0 0 loop_pad_s_7
port 26 nsew signal bidirectional
flabel metal2 267522 519384 267598 519940 0 FreeSans 1024 0 0 0 tie_pad_n_12
port 27 nsew signal bidirectional
flabel metal2 247522 518984 247598 519940 0 FreeSans 1024 0 0 0 ta_pad_n_13
port 28 nsew signal bidirectional
flabel metal2 227522 518584 227598 519940 0 FreeSans 1024 0 0 0 toe_pad_n_14
port 29 nsew signal bidirectional
flabel metal2 207522 518184 207598 519940 0 FreeSans 1024 0 0 0 ty_pad_n_15
port 30 nsew signal bidirectional
<< properties >>
string LEFclass COVER
string FIXED_BBOX 0 0 595120 595120
<< end >>
