`default_nettype none

(* blackbox *)
module tt_logo (
);

endmodule
