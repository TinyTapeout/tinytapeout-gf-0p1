magic
tech gf180mcuD
magscale 1 5
timestamp 1757269625
<< metal3 >>
rect 0 0 10028 28
<< labels >>
flabel metal3 0 0 28 28 0 FreeSans 128 0 0 0 A
port 1 nsew signal bidirectional
flabel metal3 10000 0 10028 28 0 FreeSans 128 0 0 0 B
port 2 nsew signal bidirectional
<< properties >> 
string FIXED_BBOX 0 0 10028 28
<< end >>
