magic
tech gf180mcuD
magscale 1 10
timestamp 1757387022
<< metal2 >>
rect 127240 518884 127880 520332
rect 127230 518564 127240 518884
rect 127560 518564 145880 518884
rect 145560 509872 145880 518564
rect 147240 515884 147880 520332
rect 147230 515564 147240 515884
rect 147560 510532 147880 515884
rect 147550 510212 147560 510532
rect 147880 510212 147890 510532
rect 145550 509552 145560 509872
rect 145880 509552 145890 509872
rect 138444 471720 138764 471730
rect 76236 471400 138444 471720
rect 76236 467880 76556 471400
rect 138444 471390 138764 471400
rect 74788 467240 76556 467880
rect 76236 450720 76556 467240
rect 187060 454984 188060 520444
rect 207522 518260 207598 519940
rect 227522 518660 227598 519940
rect 247522 519060 247598 519940
rect 267522 519460 267598 519940
rect 282337 519460 282413 521060
rect 267522 519384 282413 519460
rect 293940 519060 294016 521060
rect 247522 518984 294016 519060
rect 294086 518660 294162 521060
rect 227522 518584 294162 518660
rect 294232 518260 294308 521060
rect 407060 518544 408060 520444
rect 207522 518184 294308 518260
rect 401073 517544 408060 518544
rect 187050 453984 187060 454984
rect 188060 453984 188070 454984
rect 401073 453584 402073 517544
rect 427060 515544 428060 520444
rect 467240 518884 467880 520332
rect 405673 514544 428060 515544
rect 450400 518564 471720 518884
rect 405673 454984 406673 514544
rect 450400 510532 450720 518564
rect 450390 510212 450400 510532
rect 450720 510212 450730 510532
rect 471400 456332 471720 518564
rect 518564 467880 518884 467890
rect 518884 467560 520332 467880
rect 518564 467240 520332 467560
rect 471390 456012 471400 456332
rect 471720 456012 471730 456332
rect 405663 453984 405673 454984
rect 406673 453984 406683 454984
rect 401063 452584 401073 453584
rect 402073 452584 402083 453584
rect 84244 450720 84564 450730
rect 76236 450400 84244 450720
rect 84244 450390 84564 450400
rect 510000 450560 510320 450570
rect 518564 450560 518884 467240
rect 510320 450240 518884 450560
rect 510000 450230 510320 450240
rect 510660 448560 510980 448570
rect 510980 448240 512884 448560
rect 510660 448230 510980 448240
rect 512564 447560 512884 448240
rect 515564 447880 515884 447890
rect 515884 447560 520332 447880
rect 512564 447240 520332 447560
rect 74676 427060 80576 428060
rect 74676 407060 77576 408060
rect 76576 402673 77576 407060
rect 79576 406673 80576 427060
rect 454544 408060 455544 408070
rect 455544 407060 520444 408060
rect 454544 407050 455544 407060
rect 139640 406673 140640 406683
rect 79576 405673 139640 406673
rect 139640 405663 140640 405673
rect 141040 402673 142040 402683
rect 76576 401673 141040 402673
rect 141040 401663 142040 401673
rect 453144 194447 454144 194457
rect 454144 193447 518544 194447
rect 453144 193437 454144 193447
rect 454544 189447 455544 189457
rect 455544 188447 515544 189447
rect 454544 188437 455544 188447
rect 139640 188060 140640 188070
rect 74676 187060 139640 188060
rect 139640 187050 140640 187060
rect 514544 168060 515544 188447
rect 517544 188060 518544 193447
rect 517544 187060 520444 188060
rect 514544 167060 520444 168060
rect 84244 147880 84564 147890
rect 74788 147560 84244 147880
rect 74788 147240 79236 147560
rect 84244 147550 84564 147560
rect 79236 147230 79556 147240
rect 84904 145880 85224 145890
rect 76236 145560 84904 145880
rect 76236 127880 76556 145560
rect 84904 145550 85224 145560
rect 510660 143720 510980 143730
rect 510980 143400 518884 143720
rect 510660 143390 510980 143400
rect 192437 141488 192447 142488
rect 193447 141488 193457 142488
rect 188437 140088 188447 141088
rect 189447 140088 189457 141088
rect 122390 138556 122400 138876
rect 122720 138556 122730 138876
rect 74788 127560 76556 127880
rect 74788 127240 76236 127560
rect 76236 127230 76556 127240
rect 122400 76556 122720 138556
rect 145390 84244 145400 84564
rect 145720 84244 145730 84564
rect 145400 76556 145720 84244
rect 188447 80576 189447 140088
rect 122400 76236 145720 76556
rect 167060 79576 189447 80576
rect 127240 74788 127880 76236
rect 167060 74676 168060 79576
rect 192447 77576 193447 141488
rect 407050 140088 407060 141088
rect 408060 140088 408070 141088
rect 187060 76576 193447 77576
rect 187060 74676 188060 76576
rect 207522 75180 207598 76136
rect 227522 75180 227598 76136
rect 407060 74676 408060 140088
rect 518564 127880 518884 143400
rect 518564 127240 520332 127880
rect 456460 123720 456780 123730
rect 518564 123720 518884 127240
rect 456780 123400 518884 123720
rect 456460 123390 456780 123400
rect 450230 85690 450240 86010
rect 450560 85690 450570 86010
rect 448230 85030 448240 85350
rect 448560 85030 448570 85350
rect 448240 82556 448560 85030
rect 447240 82236 448560 82556
rect 447240 79236 447560 82236
rect 447880 79236 447890 79556
rect 447240 74788 447880 79236
rect 450240 76556 450560 85690
rect 450240 76236 467560 76556
rect 467880 76236 467890 76556
rect 467240 74788 467880 76236
<< via2 >>
rect 127240 518564 127560 518884
rect 147240 515564 147560 515884
rect 147560 510212 147880 510532
rect 145560 509552 145880 509872
rect 138444 471400 138764 471720
rect 187060 453984 188060 454984
rect 450400 510212 450720 510532
rect 518564 467560 518884 467880
rect 471400 456012 471720 456332
rect 405673 453984 406673 454984
rect 401073 452584 402073 453584
rect 84244 450400 84564 450720
rect 510000 450240 510320 450560
rect 510660 448240 510980 448560
rect 515564 447560 515884 447880
rect 454544 407060 455544 408060
rect 139640 405673 140640 406673
rect 141040 401673 142040 402673
rect 453144 193447 454144 194447
rect 454544 188447 455544 189447
rect 139640 187060 140640 188060
rect 84244 147560 84564 147880
rect 79236 147240 79556 147560
rect 84904 145560 85224 145880
rect 510660 143400 510980 143720
rect 192447 141488 193447 142488
rect 188447 140088 189447 141088
rect 122400 138556 122720 138876
rect 76236 127240 76556 127560
rect 145400 84244 145720 84564
rect 407060 140088 408060 141088
rect 456460 123400 456780 123720
rect 450240 85690 450560 86010
rect 448240 85030 448560 85350
rect 447560 79236 447880 79556
rect 467560 76236 467880 76556
<< metal3 >>
rect 127240 518884 127560 518894
rect 120560 518564 127240 518884
rect 120560 455448 120880 518564
rect 127240 518554 127560 518564
rect 147240 515884 147560 515894
rect 122560 515564 147240 515884
rect 122560 456108 122880 515564
rect 147240 515554 147560 515564
rect 147560 510532 147880 510541
rect 450400 510532 450720 510541
rect 147551 510212 147560 510532
rect 147880 510212 147889 510532
rect 450391 510212 450400 510532
rect 450720 510212 450729 510532
rect 147560 510203 147880 510212
rect 450400 510203 450720 510212
rect 145560 509872 145880 509881
rect 145551 509552 145560 509872
rect 145880 509552 145889 509872
rect 145560 509543 145880 509552
rect 455800 475560 456120 475570
rect 456120 475240 518884 475560
rect 455800 475230 456120 475240
rect 138444 471720 138764 471729
rect 138435 471400 138444 471720
rect 138764 471400 138773 471720
rect 456460 471560 456780 471570
rect 138444 471391 138764 471400
rect 456780 471240 515884 471560
rect 456460 471230 456780 471240
rect 471400 456332 471720 456341
rect 122550 455788 122560 456108
rect 122880 455788 122890 456108
rect 471391 456012 471400 456332
rect 471720 456012 471729 456332
rect 471400 456003 471720 456012
rect 120550 455128 120560 455448
rect 120880 455128 120890 455448
rect 187060 454984 188060 454993
rect 405673 454984 406673 454993
rect 187051 453984 187060 454984
rect 188060 453984 188069 454984
rect 405664 453984 405673 454984
rect 406673 453984 406682 454984
rect 187060 453975 188060 453984
rect 405673 453975 406673 453984
rect 401073 453584 402073 453593
rect 401064 452584 401073 453584
rect 402073 452584 402082 453584
rect 401073 452575 402073 452584
rect 84244 450720 84564 450729
rect 84235 450400 84244 450720
rect 84564 450400 84573 450720
rect 510000 450560 510320 450569
rect 84244 450391 84564 450400
rect 509991 450240 510000 450560
rect 510320 450240 510329 450560
rect 510000 450231 510320 450240
rect 510660 448560 510980 448569
rect 510651 448240 510660 448560
rect 510980 448240 510989 448560
rect 510660 448231 510980 448240
rect 515564 447880 515884 471240
rect 518564 467880 518884 475240
rect 518554 467560 518564 467880
rect 518884 467560 518894 467880
rect 515554 447560 515564 447880
rect 515884 447560 515894 447880
rect 454544 408060 455544 408069
rect 454535 407060 454544 408060
rect 455544 407060 455553 408060
rect 454544 407051 455544 407060
rect 139640 406673 140640 406682
rect 139631 405673 139640 406673
rect 140640 405673 140649 406673
rect 139640 405664 140640 405673
rect 141040 402673 142040 402682
rect 141031 401673 141040 402673
rect 142040 401673 142049 402673
rect 141040 401664 142040 401673
rect 453144 194447 454144 194456
rect 453135 193447 453144 194447
rect 454144 193447 454153 194447
rect 453144 193438 454144 193447
rect 454544 189447 455544 189456
rect 454535 188447 454544 189447
rect 455544 188447 455553 189447
rect 454544 188438 455544 188447
rect 139640 188060 140640 188069
rect 139631 187060 139640 188060
rect 140640 187060 140649 188060
rect 139640 187051 140640 187060
rect 84244 147880 84564 147889
rect 84235 147560 84244 147880
rect 84564 147560 84573 147880
rect 79226 147240 79236 147560
rect 79556 147240 79566 147560
rect 84244 147551 84564 147560
rect 76226 127240 76236 127560
rect 76556 127240 76566 127560
rect 76236 120880 76556 127240
rect 79236 122880 79556 147240
rect 84904 145880 85224 145889
rect 84895 145560 84904 145880
rect 85224 145560 85233 145880
rect 84904 145551 85224 145560
rect 510660 143720 510980 143729
rect 510651 143400 510660 143720
rect 510980 143400 510989 143720
rect 510660 143391 510980 143400
rect 192447 142488 193447 142497
rect 192438 141488 192447 142488
rect 193447 141488 193456 142488
rect 192447 141479 193447 141488
rect 188447 141088 189447 141097
rect 407060 141088 408060 141097
rect 188438 140088 188447 141088
rect 189447 140088 189456 141088
rect 407051 140088 407060 141088
rect 408060 140088 408069 141088
rect 188447 140079 189447 140088
rect 407060 140079 408060 140088
rect 474230 139400 474240 139720
rect 474560 139400 474570 139720
rect 122400 138876 122720 138885
rect 122391 138556 122400 138876
rect 122720 138556 122729 138876
rect 471230 138740 471240 139060
rect 471560 138740 471570 139060
rect 122400 138547 122720 138556
rect 456460 123720 456780 123729
rect 456451 123400 456460 123720
rect 456780 123400 456789 123720
rect 456460 123391 456780 123400
rect 138444 122880 138764 122890
rect 79236 122560 138444 122880
rect 138444 122550 138764 122560
rect 139104 120880 139424 120890
rect 76236 120560 139104 120880
rect 139104 120550 139424 120560
rect 450240 86010 450560 86019
rect 450231 85690 450240 86010
rect 450560 85690 450569 86010
rect 450240 85681 450560 85690
rect 448240 85350 448560 85359
rect 448231 85030 448240 85350
rect 448560 85030 448569 85350
rect 448240 85021 448560 85030
rect 145400 84564 145720 84573
rect 145391 84244 145400 84564
rect 145720 84244 145729 84564
rect 145400 84235 145720 84244
rect 447560 79556 447880 79566
rect 471240 79556 471560 138740
rect 447880 79236 471560 79556
rect 447560 79226 447880 79236
rect 467560 76556 467880 76566
rect 474240 76556 474560 139400
rect 467880 76236 474560 76556
rect 467560 76226 467880 76236
<< via3 >>
rect 147560 510212 147880 510532
rect 450400 510212 450720 510532
rect 145560 509552 145880 509872
rect 455800 475240 456120 475560
rect 138444 471400 138764 471720
rect 456460 471240 456780 471560
rect 122560 455788 122880 456108
rect 471400 456012 471720 456332
rect 120560 455128 120880 455448
rect 187060 453984 188060 454984
rect 405673 453984 406673 454984
rect 401073 452584 402073 453584
rect 84244 450400 84564 450720
rect 510000 450240 510320 450560
rect 510660 448240 510980 448560
rect 454544 407060 455544 408060
rect 139640 405673 140640 406673
rect 141040 401673 142040 402673
rect 453144 193447 454144 194447
rect 454544 188447 455544 189447
rect 139640 187060 140640 188060
rect 84244 147560 84564 147880
rect 84904 145560 85224 145880
rect 510660 143400 510980 143720
rect 192447 141488 193447 142488
rect 188447 140088 189447 141088
rect 407060 140088 408060 141088
rect 474240 139400 474560 139720
rect 122400 138556 122720 138876
rect 471240 138740 471560 139060
rect 456460 123400 456780 123720
rect 138444 122560 138764 122880
rect 139104 120560 139424 120880
rect 450240 85690 450560 86010
rect 448240 85030 448560 85350
rect 145400 84244 145720 84564
<< metal4 >>
rect 147560 510532 147880 510541
rect 450400 510532 450720 510541
rect 147551 510212 147560 510532
rect 147880 510212 147889 510532
rect 450391 510212 450400 510532
rect 450720 510212 450729 510532
rect 147560 510203 147880 510212
rect 450400 510203 450720 510212
rect 145560 509872 145880 509881
rect 145551 509552 145560 509872
rect 145880 509552 145889 509872
rect 145560 509543 145880 509552
rect 455800 475560 456120 476840
rect 455791 475240 455800 475560
rect 456120 475240 456129 475560
rect 138444 471720 138764 473000
rect 138435 471400 138444 471720
rect 138764 471400 138773 471720
rect 138444 470120 138764 471400
rect 455800 469960 456120 475240
rect 456460 471560 456780 476840
rect 456451 471240 456460 471560
rect 456780 471240 456789 471560
rect 456460 469960 456780 471240
rect 471400 456332 471720 456341
rect 122560 456108 122880 456117
rect 122551 455788 122560 456108
rect 122880 455788 122889 456108
rect 471391 456012 471400 456332
rect 471720 456012 471729 456332
rect 471400 456003 471720 456012
rect 122560 455779 122880 455788
rect 120560 455448 120880 455457
rect 120551 455128 120560 455448
rect 120880 455128 120889 455448
rect 120560 455119 120880 455128
rect 187060 454984 188060 454993
rect 405673 454984 406673 454993
rect 187051 453984 187060 454984
rect 188060 453984 188069 454984
rect 405664 453984 405673 454984
rect 406673 453984 406682 454984
rect 187060 453975 188060 453984
rect 405673 453975 406673 453984
rect 401073 453584 402073 453593
rect 401064 452584 401073 453584
rect 402073 452584 402082 453584
rect 401073 452575 402073 452584
rect 84244 450720 84564 452000
rect 84235 450400 84244 450720
rect 84564 450400 84573 450720
rect 510000 450560 510320 451840
rect 84244 449120 84564 450400
rect 509991 450240 510000 450560
rect 510320 450240 510329 450560
rect 510000 446960 510320 450240
rect 510660 448560 510980 451840
rect 510651 448240 510660 448560
rect 510980 448240 510989 448560
rect 510660 446960 510980 448240
rect 139640 406673 140640 410673
rect 139631 405673 139640 406673
rect 140640 405673 140649 406673
rect 139640 397673 140640 405673
rect 141040 402673 142040 410673
rect 454544 408060 455544 412060
rect 454535 407060 454544 408060
rect 455544 407060 455553 408060
rect 454544 403060 455544 407060
rect 141031 401673 141040 402673
rect 142040 401673 142049 402673
rect 141040 397673 142040 401673
rect 453144 194447 454144 198447
rect 453135 193447 453144 194447
rect 454144 193447 454153 194447
rect 139640 188060 140640 192060
rect 139631 187060 139640 188060
rect 140640 187060 140649 188060
rect 139640 183060 140640 187060
rect 453144 184447 454144 193447
rect 454544 189447 455544 198447
rect 454535 188447 454544 189447
rect 455544 188447 455553 189447
rect 454544 184447 455544 188447
rect 84244 147880 84564 149160
rect 84235 147560 84244 147880
rect 84564 147560 84573 147880
rect 84244 144280 84564 147560
rect 84904 145880 85224 149160
rect 84895 145560 84904 145880
rect 85224 145560 85233 145880
rect 84904 144280 85224 145560
rect 510660 143720 510980 145000
rect 510651 143400 510660 143720
rect 510980 143400 510989 143720
rect 192447 142488 193447 142497
rect 192438 141488 192447 142488
rect 193447 141488 193456 142488
rect 510660 142120 510980 143400
rect 192447 141479 193447 141488
rect 188447 141088 189447 141097
rect 407060 141088 408060 141097
rect 188438 140088 188447 141088
rect 189447 140088 189456 141088
rect 407051 140088 407060 141088
rect 408060 140088 408069 141088
rect 188447 140079 189447 140088
rect 407060 140079 408060 140088
rect 474240 139720 474560 139729
rect 474231 139400 474240 139720
rect 474560 139400 474569 139720
rect 474240 139391 474560 139400
rect 471240 139060 471560 139069
rect 122400 138876 122720 138885
rect 122391 138556 122400 138876
rect 122720 138556 122729 138876
rect 471231 138740 471240 139060
rect 471560 138740 471569 139060
rect 471240 138731 471560 138740
rect 122400 138547 122720 138556
rect 138444 122880 138764 124160
rect 138435 122560 138444 122880
rect 138764 122560 138773 122880
rect 138444 119280 138764 122560
rect 139104 120880 139424 124160
rect 456460 123720 456780 125000
rect 456451 123400 456460 123720
rect 456780 123400 456789 123720
rect 456460 122120 456780 123400
rect 139095 120560 139104 120880
rect 139424 120560 139433 120880
rect 139104 119280 139424 120560
rect 450240 86010 450560 86019
rect 450231 85690 450240 86010
rect 450560 85690 450569 86010
rect 450240 85681 450560 85690
rect 448240 85350 448560 85359
rect 448231 85030 448240 85350
rect 448560 85030 448569 85350
rect 448240 85021 448560 85030
rect 145400 84564 145720 84573
rect 145391 84244 145400 84564
rect 145720 84244 145729 84564
rect 145400 84235 145720 84244
<< via4 >>
rect 147560 510212 147880 510532
rect 450400 510212 450720 510532
rect 145560 509552 145880 509872
rect 122560 455788 122880 456108
rect 471400 456012 471720 456332
rect 120560 455128 120880 455448
rect 187060 453984 188060 454984
rect 405673 453984 406673 454984
rect 401073 452584 402073 453584
rect 192447 141488 193447 142488
rect 188447 140088 189447 141088
rect 407060 140088 408060 141088
rect 474240 139400 474560 139720
rect 122400 138556 122720 138876
rect 471240 138740 471560 139060
rect 450240 85690 450560 86010
rect 448240 85030 448560 85350
rect 145400 84244 145720 84564
<< metal5 >>
rect 147560 510532 147880 510541
rect 450400 510532 450720 510541
rect 144280 510212 147560 510532
rect 147880 510212 149160 510532
rect 449120 510212 450400 510532
rect 450720 510212 452000 510532
rect 147560 510203 147880 510212
rect 450400 510203 450720 510212
rect 145560 509872 145880 509881
rect 144280 509552 145560 509872
rect 145880 509552 149160 509872
rect 145560 509543 145880 509552
rect 471400 456332 471720 456341
rect 122560 456108 122880 456117
rect 119280 455788 122560 456108
rect 122880 455788 124160 456108
rect 470120 456012 471400 456332
rect 471720 456012 473000 456332
rect 471400 456003 471720 456012
rect 122560 455779 122880 455788
rect 120560 455448 120880 455457
rect 119280 455128 120560 455448
rect 120880 455128 124160 455448
rect 120560 455119 120880 455128
rect 187060 454984 188060 454993
rect 405673 454984 406673 454993
rect 183060 453984 187060 454984
rect 188060 453984 192060 454984
rect 397073 453984 405673 454984
rect 406673 453984 410673 454984
rect 187060 453975 188060 453984
rect 405673 453975 406673 453984
rect 401073 453584 402073 453593
rect 397073 452584 401073 453584
rect 402073 452584 410673 453584
rect 401073 452575 402073 452584
rect 192447 142488 193447 142497
rect 184447 141488 192447 142488
rect 193447 141488 197447 142488
rect 192447 141479 193447 141488
rect 188447 141088 189447 141097
rect 407060 141088 408060 141097
rect 184447 140088 188447 141088
rect 189447 140088 197447 141088
rect 403060 140088 407060 141088
rect 408060 140088 412060 141088
rect 188447 140079 189447 140088
rect 407060 140079 408060 140088
rect 474240 139720 474560 139729
rect 469960 139400 474240 139720
rect 474560 139400 475840 139720
rect 474240 139391 474560 139400
rect 471240 139060 471560 139069
rect 122400 138876 122720 138885
rect 121120 138556 122400 138876
rect 122720 138556 124000 138876
rect 469960 138740 471240 139060
rect 471560 138740 475840 139060
rect 471240 138731 471560 138740
rect 122400 138547 122720 138556
rect 450240 86010 450560 86019
rect 446960 85690 450240 86010
rect 450560 85690 451840 86010
rect 450240 85681 450560 85690
rect 448240 85350 448560 85359
rect 446960 85030 448240 85350
rect 448560 85030 451840 85350
rect 448240 85021 448560 85030
rect 145400 84564 145720 84573
rect 144120 84244 145400 84564
rect 145720 84244 147000 84564
rect 145400 84235 145720 84244
use power_taper  power_taper_0
timestamp 1757356513
transform 1 0 120332 0 1 74060
box 0 -200 14456 1344
use power_taper  power_taper_2
timestamp 1757356513
transform 1 0 160332 0 1 74060
box 0 -200 14456 1344
use power_taper  power_taper_3
timestamp 1757356513
transform 1 0 180332 0 1 74060
box 0 -200 14456 1344
use power_taper  power_taper_4
timestamp 1757356513
transform 1 0 400332 0 1 74060
box 0 -200 14456 1344
use power_taper  power_taper_6
timestamp 1757356513
transform 1 0 440332 0 1 74060
box 0 -200 14456 1344
use power_taper  power_taper_7
timestamp 1757356513
transform 1 0 460332 0 1 74060
box 0 -200 14456 1344
use power_taper  power_taper_8
timestamp 1757356513
transform 0 -1 521060 1 0 120332
box 0 -200 14456 1344
use power_taper  power_taper_10
timestamp 1757356513
transform 0 -1 521060 1 0 160332
box 0 -200 14456 1344
use power_taper  power_taper_11
timestamp 1757356513
transform 0 -1 521060 1 0 180332
box 0 -200 14456 1344
use power_taper  power_taper_12
timestamp 1757356513
transform 0 -1 521060 1 0 400332
box 0 -200 14456 1344
use power_taper  power_taper_14
timestamp 1757356513
transform 0 -1 521060 1 0 440332
box 0 -200 14456 1344
use power_taper  power_taper_15
timestamp 1757356513
transform 0 -1 521060 1 0 460332
box 0 -200 14456 1344
use power_taper  power_taper_16
timestamp 1757356513
transform -1 0 474788 0 -1 521060
box 0 -200 14456 1344
use power_taper  power_taper_18
timestamp 1757356513
transform -1 0 434788 0 -1 521060
box 0 -200 14456 1344
use power_taper  power_taper_19
timestamp 1757356513
transform -1 0 414788 0 -1 521060
box 0 -200 14456 1344
use power_taper  power_taper_20
timestamp 1757356513
transform -1 0 194788 0 -1 521060
box 0 -200 14456 1344
use power_taper  power_taper_22
timestamp 1757356513
transform -1 0 154788 0 -1 521060
box 0 -200 14456 1344
use power_taper  power_taper_23
timestamp 1757356513
transform -1 0 134788 0 -1 521060
box 0 -200 14456 1344
use power_taper  power_taper_24
timestamp 1757356513
transform 0 1 74060 -1 0 474788
box 0 -200 14456 1344
use power_taper  power_taper_26
timestamp 1757356513
transform 0 1 74060 -1 0 434788
box 0 -200 14456 1344
use power_taper  power_taper_27
timestamp 1757356513
transform 0 1 74060 -1 0 414788
box 0 -200 14456 1344
use power_taper  power_taper_28
timestamp 1757356513
transform 0 1 74060 -1 0 194788
box 0 -200 14456 1344
use power_taper  power_taper_30
timestamp 1757356513
transform 0 1 74060 -1 0 154788
box 0 -200 14456 1344
use power_taper  power_taper_31
timestamp 1757356513
transform 0 1 74060 -1 0 134788
box 0 -200 14456 1344
use signal_taper  signal_taper_0
timestamp 1757356446
transform 1 0 203128 0 1 74060
box 0 -200 8864 1232
use signal_taper  signal_taper_1
timestamp 1757356446
transform 1 0 223128 0 1 74060
box 0 -200 8864 1232
use signal_taper  signal_taper_2
timestamp 1757356446
transform -1 0 271992 0 -1 521060
box 0 -200 8864 1232
use signal_taper  signal_taper_3
timestamp 1757356446
transform -1 0 251992 0 -1 521060
box 0 -200 8864 1232
use signal_taper  signal_taper_4
timestamp 1757356446
transform -1 0 231992 0 -1 521060
box 0 -200 8864 1232
use signal_taper  signal_taper_5
timestamp 1757356446
transform -1 0 211992 0 -1 521060
box 0 -200 8864 1232
<< labels >>
flabel metal2 167060 74676 168060 75676 0 FreeSans 1024 0 0 0 vss_pad_s_4
port 2 nsew ground bidirectional
flabel metal2 187060 74676 188060 75676 0 FreeSans 1024 0 0 0 vddcore0_pad_s_5
port 3 nsew power bidirectional
flabel metal2 407060 74676 408060 75676 0 FreeSans 1024 0 0 0 vss_pad_s_16
port 4 nsew ground bidirectional
flabel metal2 519444 167060 520444 168060 0 FreeSans 1024 0 0 0 vss_pad_e_4
port 8 nsew ground bidirectional
flabel metal2 519444 187060 520444 188060 0 FreeSans 1024 0 0 0 vddcore0_pad_e_5
port 9 nsew power bidirectional
flabel metal2 519444 407060 520444 408060 0 FreeSans 1024 0 0 0 vss_pad_e_16
port 10 nsew ground bidirectional
flabel metal2 467240 519692 467880 520332 0 FreeSans 1024 0 0 0 vss_pad_n_2
port 13 nsew ground bidirectional
flabel metal2 427060 519444 428060 520444 0 FreeSans 1024 0 0 0 vss_pad_n_4
port 14 nsew ground bidirectional
flabel metal2 407060 519444 408060 520444 0 FreeSans 1024 0 0 0 vddcore0_pad_n_5
port 15 nsew power bidirectional
flabel metal2 187060 519444 188060 520444 0 FreeSans 1024 0 0 0 vss_pad_n_16
port 16 nsew ground bidirectional
flabel metal2 74788 467240 75428 467880 0 FreeSans 1024 0 0 0 vss_pad_w_2
port 19 nsew ground bidirectional
flabel metal2 74676 427060 75676 428060 0 FreeSans 1024 0 0 0 vss_pad_w_4
port 20 nsew ground bidirectional
flabel metal2 74676 407060 75676 408060 0 FreeSans 1024 0 0 0 vddcore0_pad_w_5
port 21 nsew power bidirectional
flabel metal2 74676 187060 75676 188060 0 FreeSans 1024 0 0 0 vss_pad_w_16
port 22 nsew ground bidirectional
flabel metal2 207522 75180 207598 76136 0 FreeSans 1024 0 0 0 loop_pad_s_6
port 25 nsew signal bidirectional
flabel metal2 227522 75180 227598 76136 0 FreeSans 1024 0 0 0 loop_pad_s_7
port 26 nsew signal bidirectional
flabel metal2 267522 519384 267598 519940 0 FreeSans 1024 0 0 0 tie_pad_n_12
port 27 nsew signal bidirectional
flabel metal2 247522 518984 247598 519940 0 FreeSans 1024 0 0 0 ta_pad_n_13
port 28 nsew signal bidirectional
flabel metal2 227522 518584 227598 519940 0 FreeSans 1024 0 0 0 toe_pad_n_14
port 29 nsew signal bidirectional
flabel metal2 207522 518184 207598 519940 0 FreeSans 1024 0 0 0 ty_pad_n_15
port 30 nsew signal bidirectional
flabel metal2 74788 147240 75428 147880 0 FreeSans 1024 0 0 0 vss_pad_w_18
port 23 nsew ground bidirectional
flabel metal2 74788 127240 75428 127880 0 FreeSans 1024 0 0 0 vddcore2_pad_w_19
port 24 nsew power bidirectional
flabel metal2 447240 74788 447880 75428 0 FreeSans 1024 0 0 0 vss_pad_s_18
port 5 nsew ground bidirectional
flabel metal2 467240 74788 467880 75428 0 FreeSans 1024 0 0 0 vddcore3_pad_s_19
port 6 nsew power bidirectional
flabel metal2 519692 447240 520332 447880 0 FreeSans 1024 0 0 0 vss_pad_e_18
port 11 nsew ground bidirectional
flabel metal2 519692 467240 520332 467880 0 FreeSans 1024 0 0 0 vddcore4_pad_e_19
port 12 nsew power bidirectional
flabel metal2 147240 519692 147880 520332 0 FreeSans 1024 0 0 0 vss_pad_n_18
port 17 nsew ground bidirectional
flabel metal2 127240 519692 127880 520332 0 FreeSans 1024 0 0 0 vddcore1_pad_n_19
port 18 nsew power bidirectional
flabel metal2 127240 74788 127880 75428 0 FreeSans 1024 0 0 0 vss_pad_s_2
port 1 nsew ground bidirectional
flabel metal2 519692 127240 520332 127880 0 FreeSans 1024 0 0 0 vss_pad_e_2
port 7 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 595120 595120
string LEFclass COVER
<< end >>
