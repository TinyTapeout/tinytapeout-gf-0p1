magic
tech gf180mcuD
magscale 1 5
timestamp 1757295381
<< metal2 >>
rect 2202 588 2230 616
rect 2201 560 2231 588
rect 2196 532 2236 560
rect 2191 504 2241 532
rect 2184 476 2248 504
rect 2174 448 2258 476
rect 2163 420 2269 448
rect 2148 392 2284 420
rect 2128 364 2304 392
rect 2104 336 2328 364
rect 2072 308 2360 336
rect 2031 280 2401 308
rect 1979 252 2453 280
rect 1912 224 2520 252
rect 1827 196 2605 224
rect 1717 168 2715 196
rect 1576 140 2856 168
rect 1396 112 3036 140
rect 1164 84 3268 112
rect 868 56 3564 84
rect 488 28 3944 56
rect 0 0 4432 28
<< end >>
