VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO loopback
  CLASS COVER ;
  FOREIGN loopback ;
  ORIGIN 0.000 0.000 ;
  SIZE 144.320 BY 44.320 ;
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 0.000 44.320 44.320 ;
    END
  END A
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 100.000 0.000 144.320 44.320 ;
    END
  END B
  OBS
      LAYER Metal2 ;
        RECT 44.320 0.000 100.000 44.320 ;
  END
END loopback
END LIBRARY

