magic
tech gf180mcuD
magscale 1 5
timestamp 1757618779
<< metal2 >>
rect 0 0 7228 800
<< end >>
