magic
tech gf180mcuD
magscale 1 5
timestamp 1757356272
<< metal2 >>
rect 136 34900 1086 35000
rect 1376 34900 2401 35000
rect 2561 34900 3586 35000
rect 3914 34900 4939 35000
rect 5099 34900 6124 35000
rect 6414 34900 7364 35000
<< end >>
