magic
tech gf180mcuD
magscale 1 10
timestamp 1757356153
<< metal2 >>
rect 3068 69800 3576 70000
rect 4204 69800 4712 70000
rect 5340 69800 5848 70000
rect 6476 69800 6984 70000
rect 8016 69800 8524 70000
rect 9152 69800 9660 70000
rect 10288 69800 10796 70000
rect 11424 69800 11932 70000
<< end >>
