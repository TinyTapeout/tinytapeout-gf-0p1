magic
tech gf180mcuD
magscale 1 10
timestamp 1757300721
<< ndiff >>
rect 147400 84904 147720 85224
<< metal2 >>
rect 207522 518260 207598 519940
rect 227522 518660 227598 519940
rect 247522 519060 247598 519940
rect 267522 519460 267598 519940
rect 282337 519460 282413 521060
rect 267522 519384 282413 519460
rect 293940 519060 294016 521060
rect 247522 518984 294016 519060
rect 294086 518660 294162 521060
rect 227522 518584 294162 518660
rect 294232 518260 294308 521060
rect 207522 518184 294308 518260
rect 188437 141488 188447 142488
rect 189447 141488 189457 142488
rect 185437 140088 185447 141088
rect 186447 140088 186457 141088
rect 147390 84904 147400 85224
rect 147720 84904 147730 85224
rect 144390 84244 144400 84564
rect 144720 84244 144730 84564
rect 144400 76556 144720 84244
rect 127400 76236 144720 76556
rect 127400 74956 127720 76236
rect 147400 74956 147720 84904
rect 185447 80576 186447 140088
rect 167060 79576 186447 80576
rect 167060 74676 168060 79576
rect 188447 77576 189447 141488
rect 187060 76576 189447 77576
rect 187060 74676 188060 76576
rect 207522 75180 207598 76136
rect 227522 75180 227598 76136
<< via2 >>
rect 188447 141488 189447 142488
rect 185447 140088 186447 141088
rect 147400 84904 147720 85224
rect 144400 84244 144720 84564
<< metal3 >>
rect 188447 142488 189447 142497
rect 188438 141488 188447 142488
rect 189447 141488 189456 142488
rect 188447 141479 189447 141488
rect 185447 141088 186447 141097
rect 185438 140088 185447 141088
rect 186447 140088 186456 141088
rect 185447 140079 186447 140088
rect 147400 85224 147720 85233
rect 147391 84904 147400 85224
rect 147720 84904 147729 85224
rect 147400 84895 147720 84904
rect 144400 84564 144720 84573
rect 144391 84244 144400 84564
rect 144720 84244 144729 84564
rect 144400 84235 144720 84244
<< via3 >>
rect 188447 141488 189447 142488
rect 185447 140088 186447 141088
rect 147400 84904 147720 85224
rect 144400 84244 144720 84564
<< metal4 >>
rect 138444 467756 138764 510532
rect 139104 468416 139424 509872
rect 180800 468416 181120 509872
rect 181460 467756 181780 510532
rect 413444 467756 413764 510532
rect 414104 468416 414424 509872
rect 455800 468416 456120 509872
rect 456460 467756 456780 510532
rect 84244 413444 84564 456108
rect 84904 414104 85224 455448
rect 87796 442634 87852 444166
rect 126600 414104 126920 455448
rect 127260 413444 127580 456108
rect 84244 138556 84564 181332
rect 84904 139216 85224 180672
rect 126600 139216 126920 180672
rect 127260 138556 127580 181332
rect 139640 140088 140640 454984
rect 141040 141488 142040 453584
rect 188447 142488 189447 142497
rect 188438 141488 188447 142488
rect 189447 141488 189456 142488
rect 453144 141488 454144 453584
rect 188447 141479 189447 141488
rect 185447 141088 186447 141097
rect 185438 140088 185447 141088
rect 186447 140088 186456 141088
rect 454544 140088 455544 454984
rect 467644 413556 467964 456332
rect 468304 414216 468624 455672
rect 510000 414216 510320 455672
rect 510660 413556 510980 456332
rect 185447 140079 186447 140088
rect 467620 138740 467940 181280
rect 468280 139400 468600 180620
rect 510000 139400 510320 180620
rect 510660 138740 510980 181280
rect 138444 84244 138764 126908
rect 139104 84904 139424 126248
rect 147400 85224 147720 85233
rect 147391 84904 147400 85224
rect 147720 84904 147729 85224
rect 180800 84904 181120 126248
rect 147400 84895 147720 84904
rect 144400 84564 144720 84573
rect 144391 84244 144400 84564
rect 144720 84244 144729 84564
rect 181460 84244 181780 126908
rect 413420 85030 413740 127490
rect 414080 85690 414400 126830
rect 455800 85690 456120 126830
rect 456460 85030 456780 127490
rect 144400 84235 144720 84244
<< via4 >>
rect 188447 141488 189447 142488
rect 185447 140088 186447 141088
rect 147400 84904 147720 85224
rect 144400 84244 144720 84564
<< metal5 >>
rect 138444 510212 181780 510532
rect 413444 510212 456780 510532
rect 139104 509552 181120 509872
rect 414104 509552 456120 509872
rect 139104 468416 181120 468736
rect 414104 468416 456120 468736
rect 138444 467756 181780 468076
rect 413444 467756 456780 468076
rect 84244 455788 127580 456108
rect 467644 456012 510980 456332
rect 84904 455128 126920 455448
rect 468304 455352 510320 455672
rect 139640 453984 455544 454984
rect 141040 452584 454144 453584
rect 84904 414104 126920 414424
rect 468304 414216 510320 414536
rect 84244 413444 127580 413764
rect 467644 413556 510980 413876
rect 84244 181012 127580 181332
rect 467620 180960 510980 181280
rect 84904 180352 126920 180672
rect 468280 180300 510320 180620
rect 188447 142488 189447 142497
rect 141040 141488 188447 142488
rect 189447 141488 454144 142488
rect 188447 141479 189447 141488
rect 185447 141088 186447 141097
rect 139640 140088 185447 141088
rect 186447 140088 455544 141088
rect 185447 140079 186447 140088
rect 84904 139216 126920 139536
rect 468280 139400 510320 139720
rect 84244 138556 127580 138876
rect 467620 138740 510980 139060
rect 413420 127170 456780 127490
rect 138444 126588 181780 126908
rect 414080 126510 456120 126830
rect 139104 125928 181120 126248
rect 414080 85690 456120 86010
rect 147400 85224 147720 85233
rect 139104 84904 147400 85224
rect 147720 84904 181120 85224
rect 413420 85030 456780 85350
rect 147400 84895 147720 84904
rect 144400 84564 144720 84573
rect 138444 84244 144400 84564
rect 144720 84244 181780 84564
rect 144400 84235 144720 84244
use power_taper  power_taper_0
timestamp 1757295289
transform 1 0 120332 0 1 74060
box 0 0 14456 1344
use power_taper  power_taper_1
timestamp 1757295289
transform 1 0 140332 0 1 74060
box 0 0 14456 1344
use power_taper  power_taper_2
timestamp 1757295289
transform 1 0 160332 0 1 74060
box 0 0 14456 1344
use power_taper  power_taper_3
timestamp 1757295289
transform 1 0 180332 0 1 74060
box 0 0 14456 1344
use power_taper  power_taper_4
timestamp 1757295289
transform 1 0 400332 0 1 74060
box 0 0 14456 1344
use power_taper  power_taper_5
timestamp 1757295289
transform 1 0 420332 0 1 74060
box 0 0 14456 1344
use power_taper  power_taper_6
timestamp 1757295289
transform 1 0 440332 0 1 74060
box 0 0 14456 1344
use power_taper  power_taper_7
timestamp 1757295289
transform 1 0 460332 0 1 74060
box 0 0 14456 1344
use power_taper  power_taper_8
timestamp 1757295289
transform 0 -1 521060 1 0 120332
box 0 0 14456 1344
use power_taper  power_taper_9
timestamp 1757295289
transform 0 -1 521060 1 0 140332
box 0 0 14456 1344
use power_taper  power_taper_10
timestamp 1757295289
transform 0 -1 521060 1 0 160332
box 0 0 14456 1344
use power_taper  power_taper_11
timestamp 1757295289
transform 0 -1 521060 1 0 180332
box 0 0 14456 1344
use power_taper  power_taper_12
timestamp 1757295289
transform 0 -1 521060 1 0 400332
box 0 0 14456 1344
use power_taper  power_taper_13
timestamp 1757295289
transform 0 -1 521060 1 0 420332
box 0 0 14456 1344
use power_taper  power_taper_14
timestamp 1757295289
transform 0 -1 521060 1 0 440332
box 0 0 14456 1344
use power_taper  power_taper_15
timestamp 1757295289
transform 0 -1 521060 1 0 460332
box 0 0 14456 1344
use power_taper  power_taper_16
timestamp 1757295289
transform -1 0 474788 0 -1 521060
box 0 0 14456 1344
use power_taper  power_taper_17
timestamp 1757295289
transform -1 0 454788 0 -1 521060
box 0 0 14456 1344
use power_taper  power_taper_18
timestamp 1757295289
transform -1 0 434788 0 -1 521060
box 0 0 14456 1344
use power_taper  power_taper_19
timestamp 1757295289
transform -1 0 414788 0 -1 521060
box 0 0 14456 1344
use power_taper  power_taper_20
timestamp 1757295289
transform -1 0 194788 0 -1 521060
box 0 0 14456 1344
use power_taper  power_taper_21
timestamp 1757295289
transform -1 0 174788 0 -1 521060
box 0 0 14456 1344
use power_taper  power_taper_22
timestamp 1757295289
transform -1 0 154788 0 -1 521060
box 0 0 14456 1344
use power_taper  power_taper_23
timestamp 1757295289
transform -1 0 134788 0 -1 521060
box 0 0 14456 1344
use power_taper  power_taper_24
timestamp 1757295289
transform 0 1 74060 -1 0 474788
box 0 0 14456 1344
use power_taper  power_taper_25
timestamp 1757295289
transform 0 1 74060 -1 0 454788
box 0 0 14456 1344
use power_taper  power_taper_26
timestamp 1757295289
transform 0 1 74060 -1 0 434788
box 0 0 14456 1344
use power_taper  power_taper_27
timestamp 1757295289
transform 0 1 74060 -1 0 414788
box 0 0 14456 1344
use power_taper  power_taper_28
timestamp 1757295289
transform 0 1 74060 -1 0 194788
box 0 0 14456 1344
use power_taper  power_taper_29
timestamp 1757295289
transform 0 1 74060 -1 0 174788
box 0 0 14456 1344
use power_taper  power_taper_30
timestamp 1757295289
transform 0 1 74060 -1 0 154788
box 0 0 14456 1344
use power_taper  power_taper_31
timestamp 1757295289
transform 0 1 74060 -1 0 134788
box 0 0 14456 1344
use signal_taper  signal_taper_0
timestamp 1757295381
transform 1 0 203128 0 1 74060
box 0 0 8864 1232
use signal_taper  signal_taper_1
timestamp 1757295381
transform 1 0 223128 0 1 74060
box 0 0 8864 1232
use signal_taper  signal_taper_2
timestamp 1757295381
transform -1 0 271992 0 -1 521060
box 0 0 8864 1232
use signal_taper  signal_taper_3
timestamp 1757295381
transform -1 0 251992 0 -1 521060
box 0 0 8864 1232
use signal_taper  signal_taper_4
timestamp 1757295381
transform -1 0 231992 0 -1 521060
box 0 0 8864 1232
use signal_taper  signal_taper_5
timestamp 1757295381
transform -1 0 211992 0 -1 521060
box 0 0 8864 1232
<< end >>
