VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wiring
  CLASS COVER ;
  FOREIGN wiring ;
  ORIGIN 0.000 0.000 ;
  SIZE 2975.600 BY 2975.600 ;
  PIN vss_pad_s_2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal2 ;
        RECT 611.950 692.780 613.650 694.380 ;
        RECT 612.000 390.780 613.600 692.780 ;
        RECT 726.950 421.220 728.650 422.820 ;
        RECT 727.000 390.780 728.600 421.220 ;
        RECT 612.000 389.180 728.600 390.780 ;
        RECT 636.200 381.940 639.400 389.180 ;
        RECT 635.970 381.660 639.630 381.940 ;
        RECT 635.450 381.380 640.150 381.660 ;
        RECT 634.790 381.100 640.810 381.380 ;
        RECT 633.940 380.820 641.660 381.100 ;
        RECT 632.850 380.540 642.750 380.820 ;
        RECT 631.450 380.260 644.150 380.540 ;
        RECT 629.660 379.980 645.940 380.260 ;
        RECT 627.370 379.700 648.230 379.980 ;
        RECT 624.420 379.420 651.180 379.700 ;
        RECT 620.650 379.140 654.950 379.420 ;
        RECT 615.810 378.860 659.790 379.140 ;
        RECT 609.610 378.580 665.990 378.860 ;
        RECT 601.660 370.300 673.940 378.580 ;
        RECT 601.660 369.300 611.160 370.300 ;
        RECT 614.060 369.300 624.310 370.300 ;
        RECT 625.910 369.300 636.160 370.300 ;
        RECT 639.440 369.300 649.690 370.300 ;
        RECT 651.290 369.300 661.540 370.300 ;
        RECT 664.440 369.300 673.940 370.300 ;
      LAYER Metal3 ;
        RECT 612.000 694.380 613.600 694.425 ;
        RECT 611.955 692.780 613.645 694.380 ;
        RECT 612.000 692.735 613.600 692.780 ;
        RECT 727.000 422.820 728.600 422.865 ;
        RECT 726.955 421.220 728.645 422.820 ;
        RECT 727.000 421.175 728.600 421.220 ;
      LAYER Metal4 ;
        RECT 612.000 694.380 613.600 694.425 ;
        RECT 611.955 692.780 613.645 694.380 ;
        RECT 612.000 692.735 613.600 692.780 ;
        RECT 727.000 422.820 728.600 422.865 ;
        RECT 726.955 421.220 728.645 422.820 ;
        RECT 727.000 421.175 728.600 421.220 ;
      LAYER Metal5 ;
        RECT 612.000 694.380 613.600 694.425 ;
        RECT 605.600 692.780 620.000 694.380 ;
        RECT 612.000 692.735 613.600 692.780 ;
        RECT 727.000 422.820 728.600 422.865 ;
        RECT 720.600 421.220 735.000 422.820 ;
        RECT 727.000 421.175 728.600 421.220 ;
    END
  END vss_pad_s_2
  PIN vss_pad_s_4
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal2 ;
        RECT 942.185 700.440 947.285 705.440 ;
        RECT 942.235 410.880 947.235 700.440 ;
        RECT 835.300 405.880 947.235 410.880 ;
        RECT 835.300 381.380 840.300 405.880 ;
        RECT 834.790 381.100 840.810 381.380 ;
        RECT 833.940 380.820 841.660 381.100 ;
        RECT 832.850 380.540 842.750 380.820 ;
        RECT 831.450 380.260 844.150 380.540 ;
        RECT 829.660 379.980 845.940 380.260 ;
        RECT 827.370 379.700 848.230 379.980 ;
        RECT 824.420 379.420 851.180 379.700 ;
        RECT 820.650 379.140 854.950 379.420 ;
        RECT 815.810 378.860 859.790 379.140 ;
        RECT 809.610 378.580 865.990 378.860 ;
        RECT 801.660 370.300 873.940 378.580 ;
        RECT 801.660 369.300 811.160 370.300 ;
        RECT 814.060 369.300 824.310 370.300 ;
        RECT 825.910 369.300 836.160 370.300 ;
        RECT 839.440 369.300 849.690 370.300 ;
        RECT 851.290 369.300 861.540 370.300 ;
        RECT 864.440 369.300 873.940 370.300 ;
      LAYER Metal3 ;
        RECT 942.235 705.440 947.235 705.485 ;
        RECT 942.190 700.440 947.280 705.440 ;
        RECT 942.235 700.395 947.235 700.440 ;
      LAYER Metal4 ;
        RECT 942.235 705.440 947.235 705.485 ;
        RECT 942.190 700.440 947.280 705.440 ;
        RECT 942.235 700.395 947.235 700.440 ;
      LAYER Metal5 ;
        RECT 942.235 705.440 947.235 705.485 ;
        RECT 922.235 700.440 987.235 705.440 ;
        RECT 942.235 700.395 947.235 700.440 ;
    END
  END vss_pad_s_4
  PIN vddcore0_pad_s_5
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal2 ;
        RECT 962.185 707.440 967.285 712.440 ;
        RECT 962.235 395.880 967.235 707.440 ;
        RECT 935.300 390.880 967.235 395.880 ;
        RECT 935.300 381.380 940.300 390.880 ;
        RECT 934.790 381.100 940.810 381.380 ;
        RECT 933.940 380.820 941.660 381.100 ;
        RECT 932.850 380.540 942.750 380.820 ;
        RECT 931.450 380.260 944.150 380.540 ;
        RECT 929.660 379.980 945.940 380.260 ;
        RECT 927.370 379.700 948.230 379.980 ;
        RECT 924.420 379.420 951.180 379.700 ;
        RECT 920.650 379.140 954.950 379.420 ;
        RECT 915.810 378.860 959.790 379.140 ;
        RECT 909.610 378.580 965.990 378.860 ;
        RECT 901.660 370.300 973.940 378.580 ;
        RECT 901.660 369.300 911.160 370.300 ;
        RECT 914.060 369.300 924.310 370.300 ;
        RECT 925.910 369.300 936.160 370.300 ;
        RECT 939.440 369.300 949.690 370.300 ;
        RECT 951.290 369.300 961.540 370.300 ;
        RECT 964.440 369.300 973.940 370.300 ;
      LAYER Metal3 ;
        RECT 962.235 712.440 967.235 712.485 ;
        RECT 962.190 707.440 967.280 712.440 ;
        RECT 962.235 707.395 967.235 707.440 ;
      LAYER Metal4 ;
        RECT 962.235 712.440 967.235 712.485 ;
        RECT 962.190 707.440 967.280 712.440 ;
        RECT 962.235 707.395 967.235 707.440 ;
      LAYER Metal5 ;
        RECT 962.235 712.440 967.235 712.485 ;
        RECT 922.235 707.440 987.235 712.440 ;
        RECT 962.235 707.395 967.235 707.440 ;
    END
  END vddcore0_pad_s_5
  PIN vss_pad_s_16
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal2 ;
        RECT 2035.250 700.440 2040.350 705.440 ;
        RECT 2035.300 381.380 2040.300 700.440 ;
        RECT 2034.790 381.100 2040.810 381.380 ;
        RECT 2033.940 380.820 2041.660 381.100 ;
        RECT 2032.850 380.540 2042.750 380.820 ;
        RECT 2031.450 380.260 2044.150 380.540 ;
        RECT 2029.660 379.980 2045.940 380.260 ;
        RECT 2027.370 379.700 2048.230 379.980 ;
        RECT 2024.420 379.420 2051.180 379.700 ;
        RECT 2020.650 379.140 2054.950 379.420 ;
        RECT 2015.810 378.860 2059.790 379.140 ;
        RECT 2009.610 378.580 2065.990 378.860 ;
        RECT 2001.660 370.300 2073.940 378.580 ;
        RECT 2001.660 369.300 2011.160 370.300 ;
        RECT 2014.060 369.300 2024.310 370.300 ;
        RECT 2025.910 369.300 2036.160 370.300 ;
        RECT 2039.440 369.300 2049.690 370.300 ;
        RECT 2051.290 369.300 2061.540 370.300 ;
        RECT 2064.440 369.300 2073.940 370.300 ;
      LAYER Metal3 ;
        RECT 2035.300 705.440 2040.300 705.485 ;
        RECT 2035.255 700.440 2040.345 705.440 ;
        RECT 2035.300 700.395 2040.300 700.440 ;
      LAYER Metal4 ;
        RECT 2035.300 705.440 2040.300 705.485 ;
        RECT 2035.255 700.440 2040.345 705.440 ;
        RECT 2035.300 700.395 2040.300 700.440 ;
      LAYER Metal5 ;
        RECT 2035.300 705.440 2040.300 705.485 ;
        RECT 2015.300 700.440 2060.300 705.440 ;
        RECT 2035.300 700.395 2040.300 700.440 ;
    END
  END vss_pad_s_16
  PIN vss_pad_s_18
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal2 ;
        RECT 2241.150 425.150 2242.850 426.750 ;
        RECT 2241.200 412.780 2242.800 425.150 ;
        RECT 2236.200 411.180 2242.800 412.780 ;
        RECT 2236.200 401.780 2237.800 411.180 ;
        RECT 2236.200 400.180 2239.450 401.780 ;
        RECT 2236.200 381.940 2239.400 400.180 ;
        RECT 2235.970 381.660 2239.630 381.940 ;
        RECT 2235.450 381.380 2240.150 381.660 ;
        RECT 2234.790 381.100 2240.810 381.380 ;
        RECT 2233.940 380.820 2241.660 381.100 ;
        RECT 2232.850 380.540 2242.750 380.820 ;
        RECT 2231.450 380.260 2244.150 380.540 ;
        RECT 2229.660 379.980 2245.940 380.260 ;
        RECT 2227.370 379.700 2248.230 379.980 ;
        RECT 2224.420 379.420 2251.180 379.700 ;
        RECT 2220.650 379.140 2254.950 379.420 ;
        RECT 2215.810 378.860 2259.790 379.140 ;
        RECT 2209.610 378.580 2265.990 378.860 ;
        RECT 2201.660 370.300 2273.940 378.580 ;
        RECT 2201.660 369.300 2211.160 370.300 ;
        RECT 2214.060 369.300 2224.310 370.300 ;
        RECT 2225.910 369.300 2236.160 370.300 ;
        RECT 2239.440 369.300 2249.690 370.300 ;
        RECT 2251.290 369.300 2261.540 370.300 ;
        RECT 2264.440 369.300 2273.940 370.300 ;
      LAYER Metal3 ;
        RECT 2356.150 693.700 2357.850 695.300 ;
        RECT 2241.200 426.750 2242.800 426.795 ;
        RECT 2241.155 425.150 2242.845 426.750 ;
        RECT 2241.200 425.105 2242.800 425.150 ;
        RECT 2237.800 401.780 2239.400 401.830 ;
        RECT 2356.200 401.780 2357.800 693.700 ;
        RECT 2237.800 400.180 2357.800 401.780 ;
        RECT 2237.800 400.130 2239.400 400.180 ;
      LAYER Metal4 ;
        RECT 2356.200 695.300 2357.800 695.345 ;
        RECT 2356.155 693.700 2357.845 695.300 ;
        RECT 2356.200 693.655 2357.800 693.700 ;
        RECT 2241.200 426.750 2242.800 426.795 ;
        RECT 2241.155 425.150 2242.845 426.750 ;
        RECT 2241.200 425.105 2242.800 425.150 ;
      LAYER Metal5 ;
        RECT 2356.200 695.300 2357.800 695.345 ;
        RECT 2349.800 693.700 2379.200 695.300 ;
        RECT 2356.200 693.655 2357.800 693.700 ;
        RECT 2241.200 426.750 2242.800 426.795 ;
        RECT 2234.800 425.150 2259.200 426.750 ;
        RECT 2241.200 425.105 2242.800 425.150 ;
    END
  END vss_pad_s_18
  PIN vddcore3_pad_s_19
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal2 ;
        RECT 2251.150 428.450 2252.850 430.050 ;
        RECT 2251.200 390.780 2252.800 428.450 ;
        RECT 2251.200 389.180 2339.450 390.780 ;
        RECT 2336.200 381.940 2339.400 389.180 ;
        RECT 2335.970 381.660 2339.630 381.940 ;
        RECT 2335.450 381.380 2340.150 381.660 ;
        RECT 2334.790 381.100 2340.810 381.380 ;
        RECT 2333.940 380.820 2341.660 381.100 ;
        RECT 2332.850 380.540 2342.750 380.820 ;
        RECT 2331.450 380.260 2344.150 380.540 ;
        RECT 2329.660 379.980 2345.940 380.260 ;
        RECT 2327.370 379.700 2348.230 379.980 ;
        RECT 2324.420 379.420 2351.180 379.700 ;
        RECT 2320.650 379.140 2354.950 379.420 ;
        RECT 2315.810 378.860 2359.790 379.140 ;
        RECT 2309.610 378.580 2365.990 378.860 ;
        RECT 2301.660 370.300 2373.940 378.580 ;
        RECT 2301.660 369.300 2311.160 370.300 ;
        RECT 2314.060 369.300 2324.310 370.300 ;
        RECT 2325.910 369.300 2336.160 370.300 ;
        RECT 2339.440 369.300 2349.690 370.300 ;
        RECT 2351.290 369.300 2361.540 370.300 ;
        RECT 2364.440 369.300 2373.940 370.300 ;
      LAYER Metal3 ;
        RECT 2371.150 697.000 2372.850 698.600 ;
        RECT 2251.200 430.050 2252.800 430.095 ;
        RECT 2251.155 428.450 2252.845 430.050 ;
        RECT 2251.200 428.405 2252.800 428.450 ;
        RECT 2337.800 390.780 2339.400 390.830 ;
        RECT 2371.200 390.780 2372.800 697.000 ;
        RECT 2337.800 389.180 2372.800 390.780 ;
        RECT 2337.800 389.130 2339.400 389.180 ;
      LAYER Metal4 ;
        RECT 2371.200 698.600 2372.800 698.645 ;
        RECT 2371.155 697.000 2372.845 698.600 ;
        RECT 2371.200 696.955 2372.800 697.000 ;
        RECT 2251.200 430.050 2252.800 430.095 ;
        RECT 2251.155 428.450 2252.845 430.050 ;
        RECT 2251.200 428.405 2252.800 428.450 ;
      LAYER Metal5 ;
        RECT 2371.200 698.600 2372.800 698.645 ;
        RECT 2349.800 697.000 2379.200 698.600 ;
        RECT 2371.200 696.955 2372.800 697.000 ;
        RECT 2251.200 430.050 2252.800 430.095 ;
        RECT 2234.800 428.450 2259.200 430.050 ;
        RECT 2251.200 428.405 2252.800 428.450 ;
    END
  END vddcore3_pad_s_19
  PIN vss_pad_e_2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal2 ;
        RECT 2553.300 718.600 2554.900 718.650 ;
        RECT 2553.300 717.000 2586.420 718.600 ;
        RECT 2553.300 716.950 2554.900 717.000 ;
        RECT 2584.820 639.400 2586.420 717.000 ;
        RECT 2597.020 665.990 2606.300 673.940 ;
        RECT 2596.740 664.440 2606.300 665.990 ;
        RECT 2596.740 661.540 2605.300 664.440 ;
        RECT 2596.740 659.790 2606.300 661.540 ;
        RECT 2596.460 654.950 2606.300 659.790 ;
        RECT 2596.180 651.290 2606.300 654.950 ;
        RECT 2596.180 651.180 2605.300 651.290 ;
        RECT 2595.900 649.690 2605.300 651.180 ;
        RECT 2595.900 648.230 2606.300 649.690 ;
        RECT 2595.620 645.940 2606.300 648.230 ;
        RECT 2595.340 644.150 2606.300 645.940 ;
        RECT 2595.060 642.750 2606.300 644.150 ;
        RECT 2594.780 641.660 2606.300 642.750 ;
        RECT 2594.500 640.810 2606.300 641.660 ;
        RECT 2594.220 640.150 2606.300 640.810 ;
        RECT 2593.940 639.630 2606.300 640.150 ;
        RECT 2593.660 639.440 2606.300 639.630 ;
        RECT 2593.660 639.400 2605.300 639.440 ;
        RECT 2584.820 636.200 2605.300 639.400 ;
        RECT 2282.300 618.600 2283.900 618.650 ;
        RECT 2584.820 618.600 2586.420 636.200 ;
        RECT 2593.660 636.160 2605.300 636.200 ;
        RECT 2593.660 635.970 2606.300 636.160 ;
        RECT 2593.940 635.450 2606.300 635.970 ;
        RECT 2594.220 634.790 2606.300 635.450 ;
        RECT 2594.500 633.940 2606.300 634.790 ;
        RECT 2594.780 632.850 2606.300 633.940 ;
        RECT 2595.060 631.450 2606.300 632.850 ;
        RECT 2595.340 629.660 2606.300 631.450 ;
        RECT 2595.620 627.370 2606.300 629.660 ;
        RECT 2595.900 625.910 2606.300 627.370 ;
        RECT 2595.900 624.420 2605.300 625.910 ;
        RECT 2596.180 624.310 2605.300 624.420 ;
        RECT 2596.180 620.650 2606.300 624.310 ;
        RECT 2282.300 617.000 2586.420 618.600 ;
        RECT 2282.300 616.950 2283.900 617.000 ;
        RECT 2596.460 615.810 2606.300 620.650 ;
        RECT 2596.740 614.060 2606.300 615.810 ;
        RECT 2596.740 611.160 2605.300 614.060 ;
        RECT 2596.740 609.610 2606.300 611.160 ;
        RECT 2597.020 601.660 2606.300 609.610 ;
      LAYER Metal3 ;
        RECT 2553.300 718.600 2554.900 718.645 ;
        RECT 2553.255 717.000 2554.945 718.600 ;
        RECT 2553.300 716.955 2554.900 717.000 ;
        RECT 2282.300 618.600 2283.900 618.645 ;
        RECT 2282.255 617.000 2283.945 618.600 ;
        RECT 2282.300 616.955 2283.900 617.000 ;
      LAYER Metal4 ;
        RECT 2553.300 718.600 2554.900 725.000 ;
        RECT 2553.255 717.000 2554.945 718.600 ;
        RECT 2553.300 710.600 2554.900 717.000 ;
        RECT 2282.300 618.600 2283.900 625.000 ;
        RECT 2282.255 617.000 2283.945 618.600 ;
        RECT 2282.300 610.600 2283.900 617.000 ;
    END
  END vss_pad_e_2
  PIN vss_pad_e_4
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal2 ;
        RECT 2272.720 947.235 2277.720 947.285 ;
        RECT 2272.720 942.235 2569.720 947.235 ;
        RECT 2272.720 942.185 2277.720 942.235 ;
        RECT 2564.720 840.300 2569.720 942.235 ;
        RECT 2597.020 865.990 2606.300 873.940 ;
        RECT 2596.740 864.440 2606.300 865.990 ;
        RECT 2596.740 861.540 2605.300 864.440 ;
        RECT 2596.740 859.790 2606.300 861.540 ;
        RECT 2596.460 854.950 2606.300 859.790 ;
        RECT 2596.180 851.290 2606.300 854.950 ;
        RECT 2596.180 851.180 2605.300 851.290 ;
        RECT 2595.900 849.690 2605.300 851.180 ;
        RECT 2595.900 848.230 2606.300 849.690 ;
        RECT 2595.620 845.940 2606.300 848.230 ;
        RECT 2595.340 844.150 2606.300 845.940 ;
        RECT 2595.060 842.750 2606.300 844.150 ;
        RECT 2594.780 841.660 2606.300 842.750 ;
        RECT 2594.500 840.810 2606.300 841.660 ;
        RECT 2594.220 840.300 2606.300 840.810 ;
        RECT 2564.720 839.440 2606.300 840.300 ;
        RECT 2564.720 836.160 2605.300 839.440 ;
        RECT 2564.720 835.300 2606.300 836.160 ;
        RECT 2594.220 834.790 2606.300 835.300 ;
        RECT 2594.500 833.940 2606.300 834.790 ;
        RECT 2594.780 832.850 2606.300 833.940 ;
        RECT 2595.060 831.450 2606.300 832.850 ;
        RECT 2595.340 829.660 2606.300 831.450 ;
        RECT 2595.620 827.370 2606.300 829.660 ;
        RECT 2595.900 825.910 2606.300 827.370 ;
        RECT 2595.900 824.420 2605.300 825.910 ;
        RECT 2596.180 824.310 2605.300 824.420 ;
        RECT 2596.180 820.650 2606.300 824.310 ;
        RECT 2596.460 815.810 2606.300 820.650 ;
        RECT 2596.740 814.060 2606.300 815.810 ;
        RECT 2596.740 811.160 2605.300 814.060 ;
        RECT 2596.740 809.610 2606.300 811.160 ;
        RECT 2597.020 801.660 2606.300 809.610 ;
      LAYER Metal3 ;
        RECT 2272.720 947.235 2277.720 947.280 ;
        RECT 2272.675 942.235 2277.765 947.235 ;
        RECT 2272.720 942.190 2277.720 942.235 ;
      LAYER Metal4 ;
        RECT 2272.720 947.235 2277.720 992.235 ;
        RECT 2272.675 942.235 2277.765 947.235 ;
        RECT 2272.720 922.235 2277.720 942.235 ;
    END
  END vss_pad_e_4
  PIN vddcore0_pad_e_5
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal2 ;
        RECT 2265.720 972.235 2270.720 972.285 ;
        RECT 2265.720 967.235 2584.720 972.235 ;
        RECT 2265.720 967.185 2270.720 967.235 ;
        RECT 2579.720 940.300 2584.720 967.235 ;
        RECT 2597.020 965.990 2606.300 973.940 ;
        RECT 2596.740 964.440 2606.300 965.990 ;
        RECT 2596.740 961.540 2605.300 964.440 ;
        RECT 2596.740 959.790 2606.300 961.540 ;
        RECT 2596.460 954.950 2606.300 959.790 ;
        RECT 2596.180 951.290 2606.300 954.950 ;
        RECT 2596.180 951.180 2605.300 951.290 ;
        RECT 2595.900 949.690 2605.300 951.180 ;
        RECT 2595.900 948.230 2606.300 949.690 ;
        RECT 2595.620 945.940 2606.300 948.230 ;
        RECT 2595.340 944.150 2606.300 945.940 ;
        RECT 2595.060 942.750 2606.300 944.150 ;
        RECT 2594.780 941.660 2606.300 942.750 ;
        RECT 2594.500 940.810 2606.300 941.660 ;
        RECT 2594.220 940.300 2606.300 940.810 ;
        RECT 2579.720 939.440 2606.300 940.300 ;
        RECT 2579.720 936.160 2605.300 939.440 ;
        RECT 2579.720 935.300 2606.300 936.160 ;
        RECT 2594.220 934.790 2606.300 935.300 ;
        RECT 2594.500 933.940 2606.300 934.790 ;
        RECT 2594.780 932.850 2606.300 933.940 ;
        RECT 2595.060 931.450 2606.300 932.850 ;
        RECT 2595.340 929.660 2606.300 931.450 ;
        RECT 2595.620 927.370 2606.300 929.660 ;
        RECT 2595.900 925.910 2606.300 927.370 ;
        RECT 2595.900 924.420 2605.300 925.910 ;
        RECT 2596.180 924.310 2605.300 924.420 ;
        RECT 2596.180 920.650 2606.300 924.310 ;
        RECT 2596.460 915.810 2606.300 920.650 ;
        RECT 2596.740 914.060 2606.300 915.810 ;
        RECT 2596.740 911.160 2605.300 914.060 ;
        RECT 2596.740 909.610 2606.300 911.160 ;
        RECT 2597.020 901.660 2606.300 909.610 ;
      LAYER Metal3 ;
        RECT 2265.720 972.235 2270.720 972.280 ;
        RECT 2265.675 967.235 2270.765 972.235 ;
        RECT 2265.720 967.190 2270.720 967.235 ;
      LAYER Metal4 ;
        RECT 2265.720 972.235 2270.720 992.235 ;
        RECT 2265.675 967.235 2270.765 972.235 ;
        RECT 2265.720 922.235 2270.720 967.235 ;
    END
  END vddcore0_pad_e_5
  PIN vss_pad_e_16
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal2 ;
        RECT 2597.020 2065.990 2606.300 2073.940 ;
        RECT 2596.740 2064.440 2606.300 2065.990 ;
        RECT 2596.740 2061.540 2605.300 2064.440 ;
        RECT 2596.740 2059.790 2606.300 2061.540 ;
        RECT 2596.460 2054.950 2606.300 2059.790 ;
        RECT 2596.180 2051.290 2606.300 2054.950 ;
        RECT 2596.180 2051.180 2605.300 2051.290 ;
        RECT 2595.900 2049.690 2605.300 2051.180 ;
        RECT 2595.900 2048.230 2606.300 2049.690 ;
        RECT 2595.620 2045.940 2606.300 2048.230 ;
        RECT 2595.340 2044.150 2606.300 2045.940 ;
        RECT 2595.060 2042.750 2606.300 2044.150 ;
        RECT 2594.780 2041.660 2606.300 2042.750 ;
        RECT 2594.500 2040.810 2606.300 2041.660 ;
        RECT 2272.720 2040.300 2277.720 2040.350 ;
        RECT 2594.220 2040.300 2606.300 2040.810 ;
        RECT 2272.720 2039.440 2606.300 2040.300 ;
        RECT 2272.720 2036.160 2605.300 2039.440 ;
        RECT 2272.720 2035.300 2606.300 2036.160 ;
        RECT 2272.720 2035.250 2277.720 2035.300 ;
        RECT 2594.220 2034.790 2606.300 2035.300 ;
        RECT 2594.500 2033.940 2606.300 2034.790 ;
        RECT 2594.780 2032.850 2606.300 2033.940 ;
        RECT 2595.060 2031.450 2606.300 2032.850 ;
        RECT 2595.340 2029.660 2606.300 2031.450 ;
        RECT 2595.620 2027.370 2606.300 2029.660 ;
        RECT 2595.900 2025.910 2606.300 2027.370 ;
        RECT 2595.900 2024.420 2605.300 2025.910 ;
        RECT 2596.180 2024.310 2605.300 2024.420 ;
        RECT 2596.180 2020.650 2606.300 2024.310 ;
        RECT 2596.460 2015.810 2606.300 2020.650 ;
        RECT 2596.740 2014.060 2606.300 2015.810 ;
        RECT 2596.740 2011.160 2605.300 2014.060 ;
        RECT 2596.740 2009.610 2606.300 2011.160 ;
        RECT 2597.020 2001.660 2606.300 2009.610 ;
      LAYER Metal3 ;
        RECT 2272.720 2040.300 2277.720 2040.345 ;
        RECT 2272.675 2035.300 2277.765 2040.300 ;
        RECT 2272.720 2035.255 2277.720 2035.300 ;
      LAYER Metal4 ;
        RECT 2272.720 2040.300 2277.720 2060.300 ;
        RECT 2272.675 2035.300 2277.765 2040.300 ;
        RECT 2272.720 2015.300 2277.720 2035.300 ;
    END
  END vss_pad_e_16
  PIN vss_pad_e_18
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal2 ;
        RECT 2597.020 2265.990 2606.300 2273.940 ;
        RECT 2596.740 2264.440 2606.300 2265.990 ;
        RECT 2596.740 2261.540 2605.300 2264.440 ;
        RECT 2596.740 2259.790 2606.300 2261.540 ;
        RECT 2596.460 2254.950 2606.300 2259.790 ;
        RECT 2596.180 2251.290 2606.300 2254.950 ;
        RECT 2596.180 2251.180 2605.300 2251.290 ;
        RECT 2595.900 2249.690 2605.300 2251.180 ;
        RECT 2595.900 2248.230 2606.300 2249.690 ;
        RECT 2595.620 2245.940 2606.300 2248.230 ;
        RECT 2595.340 2244.150 2606.300 2245.940 ;
        RECT 2553.300 2242.800 2554.900 2242.850 ;
        RECT 2553.300 2241.200 2564.420 2242.800 ;
        RECT 2595.060 2242.750 2606.300 2244.150 ;
        RECT 2594.780 2241.660 2606.300 2242.750 ;
        RECT 2553.300 2241.150 2554.900 2241.200 ;
        RECT 2562.820 2237.800 2564.420 2241.200 ;
        RECT 2594.500 2240.810 2606.300 2241.660 ;
        RECT 2594.220 2240.150 2606.300 2240.810 ;
        RECT 2593.940 2239.630 2606.300 2240.150 ;
        RECT 2573.820 2239.400 2575.420 2239.450 ;
        RECT 2593.660 2239.440 2606.300 2239.630 ;
        RECT 2593.660 2239.400 2605.300 2239.440 ;
        RECT 2573.820 2237.800 2605.300 2239.400 ;
        RECT 2562.820 2236.200 2605.300 2237.800 ;
        RECT 2593.660 2236.160 2605.300 2236.200 ;
        RECT 2593.660 2235.970 2606.300 2236.160 ;
        RECT 2593.940 2235.450 2606.300 2235.970 ;
        RECT 2594.220 2234.790 2606.300 2235.450 ;
        RECT 2594.500 2233.940 2606.300 2234.790 ;
        RECT 2594.780 2232.850 2606.300 2233.940 ;
        RECT 2595.060 2231.450 2606.300 2232.850 ;
        RECT 2595.340 2229.660 2606.300 2231.450 ;
        RECT 2595.620 2227.370 2606.300 2229.660 ;
        RECT 2595.900 2225.910 2606.300 2227.370 ;
        RECT 2595.900 2224.420 2605.300 2225.910 ;
        RECT 2596.180 2224.310 2605.300 2224.420 ;
        RECT 2596.180 2220.650 2606.300 2224.310 ;
        RECT 2596.460 2215.810 2606.300 2220.650 ;
        RECT 2596.740 2214.060 2606.300 2215.810 ;
        RECT 2596.740 2211.160 2605.300 2214.060 ;
        RECT 2596.740 2209.610 2606.300 2211.160 ;
        RECT 2597.020 2201.660 2606.300 2209.610 ;
      LAYER Metal3 ;
        RECT 2282.300 2357.800 2283.900 2357.850 ;
        RECT 2282.300 2356.200 2575.420 2357.800 ;
        RECT 2282.300 2356.150 2283.900 2356.200 ;
        RECT 2553.300 2242.800 2554.900 2242.845 ;
        RECT 2553.255 2241.200 2554.945 2242.800 ;
        RECT 2553.300 2241.155 2554.900 2241.200 ;
        RECT 2573.820 2239.400 2575.420 2356.200 ;
        RECT 2573.770 2237.800 2575.470 2239.400 ;
      LAYER Metal4 ;
        RECT 2282.300 2357.800 2283.900 2385.800 ;
        RECT 2282.255 2356.200 2283.945 2357.800 ;
        RECT 2282.300 2349.800 2283.900 2356.200 ;
        RECT 2553.300 2242.800 2554.900 2259.200 ;
        RECT 2553.255 2241.200 2554.945 2242.800 ;
        RECT 2553.300 2234.800 2554.900 2241.200 ;
    END
  END vss_pad_e_18
  PIN vddcore4_pad_e_19
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal2 ;
        RECT 2597.020 2365.990 2606.300 2373.940 ;
        RECT 2596.740 2364.440 2606.300 2365.990 ;
        RECT 2596.740 2361.540 2605.300 2364.440 ;
        RECT 2596.740 2359.790 2606.300 2361.540 ;
        RECT 2596.460 2354.950 2606.300 2359.790 ;
        RECT 2596.180 2351.290 2606.300 2354.950 ;
        RECT 2596.180 2351.180 2605.300 2351.290 ;
        RECT 2595.900 2349.690 2605.300 2351.180 ;
        RECT 2595.900 2348.230 2606.300 2349.690 ;
        RECT 2595.620 2345.940 2606.300 2348.230 ;
        RECT 2595.340 2344.150 2606.300 2345.940 ;
        RECT 2595.060 2342.750 2606.300 2344.150 ;
        RECT 2594.780 2341.660 2606.300 2342.750 ;
        RECT 2594.500 2340.810 2606.300 2341.660 ;
        RECT 2594.220 2340.150 2606.300 2340.810 ;
        RECT 2593.940 2339.630 2606.300 2340.150 ;
        RECT 2584.820 2339.400 2586.420 2339.450 ;
        RECT 2593.660 2339.440 2606.300 2339.630 ;
        RECT 2593.660 2339.400 2605.300 2339.440 ;
        RECT 2584.820 2336.200 2605.300 2339.400 ;
        RECT 2550.000 2252.800 2551.600 2252.850 ;
        RECT 2584.820 2252.800 2586.420 2336.200 ;
        RECT 2593.660 2336.160 2605.300 2336.200 ;
        RECT 2593.660 2335.970 2606.300 2336.160 ;
        RECT 2593.940 2335.450 2606.300 2335.970 ;
        RECT 2594.220 2334.790 2606.300 2335.450 ;
        RECT 2594.500 2333.940 2606.300 2334.790 ;
        RECT 2594.780 2332.850 2606.300 2333.940 ;
        RECT 2595.060 2331.450 2606.300 2332.850 ;
        RECT 2595.340 2329.660 2606.300 2331.450 ;
        RECT 2595.620 2327.370 2606.300 2329.660 ;
        RECT 2595.900 2325.910 2606.300 2327.370 ;
        RECT 2595.900 2324.420 2605.300 2325.910 ;
        RECT 2596.180 2324.310 2605.300 2324.420 ;
        RECT 2596.180 2320.650 2606.300 2324.310 ;
        RECT 2596.460 2315.810 2606.300 2320.650 ;
        RECT 2596.740 2314.060 2606.300 2315.810 ;
        RECT 2596.740 2311.160 2605.300 2314.060 ;
        RECT 2596.740 2309.610 2606.300 2311.160 ;
        RECT 2597.020 2301.660 2606.300 2309.610 ;
        RECT 2550.000 2251.200 2586.420 2252.800 ;
        RECT 2550.000 2251.150 2551.600 2251.200 ;
      LAYER Metal3 ;
        RECT 2279.000 2379.400 2280.600 2379.450 ;
        RECT 2279.000 2377.800 2298.900 2379.400 ;
        RECT 2279.000 2377.750 2280.600 2377.800 ;
        RECT 2297.300 2376.200 2586.420 2377.800 ;
        RECT 2584.820 2339.400 2586.420 2376.200 ;
        RECT 2584.770 2337.800 2586.470 2339.400 ;
        RECT 2550.000 2252.800 2551.600 2252.845 ;
        RECT 2549.955 2251.200 2551.645 2252.800 ;
        RECT 2550.000 2251.155 2551.600 2251.200 ;
      LAYER Metal4 ;
        RECT 2279.000 2379.400 2280.600 2385.800 ;
        RECT 2278.955 2377.800 2280.645 2379.400 ;
        RECT 2279.000 2349.800 2280.600 2377.800 ;
        RECT 2550.000 2252.800 2551.600 2259.200 ;
        RECT 2549.955 2251.200 2551.645 2252.800 ;
        RECT 2550.000 2234.800 2551.600 2251.200 ;
    END
  END vddcore4_pad_e_19
  PIN vss_pad_n_2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal2 ;
        RECT 2301.660 2605.300 2311.160 2606.300 ;
        RECT 2314.060 2605.300 2324.310 2606.300 ;
        RECT 2325.910 2605.300 2336.160 2606.300 ;
        RECT 2339.440 2605.300 2349.690 2606.300 ;
        RECT 2351.290 2605.300 2361.540 2606.300 ;
        RECT 2364.440 2605.300 2373.940 2606.300 ;
        RECT 2301.660 2597.020 2373.940 2605.300 ;
        RECT 2309.610 2596.740 2365.990 2597.020 ;
        RECT 2315.810 2596.460 2359.790 2596.740 ;
        RECT 2320.650 2596.180 2354.950 2596.460 ;
        RECT 2324.420 2595.900 2351.180 2596.180 ;
        RECT 2327.370 2595.620 2348.230 2595.900 ;
        RECT 2329.660 2595.340 2345.940 2595.620 ;
        RECT 2331.450 2595.060 2344.150 2595.340 ;
        RECT 2332.850 2594.780 2342.750 2595.060 ;
        RECT 2333.940 2594.500 2341.660 2594.780 ;
        RECT 2334.790 2594.220 2340.810 2594.500 ;
        RECT 2335.450 2593.940 2340.150 2594.220 ;
        RECT 2335.970 2593.660 2339.630 2593.940 ;
        RECT 2336.200 2586.420 2339.400 2593.660 ;
        RECT 2252.000 2584.820 2358.600 2586.420 ;
        RECT 2252.000 2552.660 2253.600 2584.820 ;
        RECT 2251.950 2551.060 2253.650 2552.660 ;
        RECT 2357.000 2281.660 2358.600 2584.820 ;
        RECT 2356.950 2280.060 2358.650 2281.660 ;
      LAYER Metal3 ;
        RECT 2252.000 2552.660 2253.600 2552.705 ;
        RECT 2251.955 2551.060 2253.645 2552.660 ;
        RECT 2252.000 2551.015 2253.600 2551.060 ;
        RECT 2357.000 2281.660 2358.600 2281.705 ;
        RECT 2356.955 2280.060 2358.645 2281.660 ;
        RECT 2357.000 2280.015 2358.600 2280.060 ;
      LAYER Metal4 ;
        RECT 2252.000 2552.660 2253.600 2552.705 ;
        RECT 2251.955 2551.060 2253.645 2552.660 ;
        RECT 2252.000 2551.015 2253.600 2551.060 ;
        RECT 2357.000 2281.660 2358.600 2281.705 ;
        RECT 2356.955 2280.060 2358.645 2281.660 ;
        RECT 2357.000 2280.015 2358.600 2280.060 ;
      LAYER Metal5 ;
        RECT 2252.000 2552.660 2253.600 2552.705 ;
        RECT 2245.600 2551.060 2260.000 2552.660 ;
        RECT 2252.000 2551.015 2253.600 2551.060 ;
        RECT 2357.000 2281.660 2358.600 2281.705 ;
        RECT 2350.600 2280.060 2365.000 2281.660 ;
        RECT 2357.000 2280.015 2358.600 2280.060 ;
    END
  END vss_pad_n_2
  PIN vss_pad_n_4
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal2 ;
        RECT 2101.660 2605.300 2111.160 2606.300 ;
        RECT 2114.060 2605.300 2124.310 2606.300 ;
        RECT 2125.910 2605.300 2136.160 2606.300 ;
        RECT 2139.440 2605.300 2149.690 2606.300 ;
        RECT 2151.290 2605.300 2161.540 2606.300 ;
        RECT 2164.440 2605.300 2173.940 2606.300 ;
        RECT 2101.660 2597.020 2173.940 2605.300 ;
        RECT 2109.610 2596.740 2165.990 2597.020 ;
        RECT 2115.810 2596.460 2159.790 2596.740 ;
        RECT 2120.650 2596.180 2154.950 2596.460 ;
        RECT 2124.420 2595.900 2151.180 2596.180 ;
        RECT 2127.370 2595.620 2148.230 2595.900 ;
        RECT 2129.660 2595.340 2145.940 2595.620 ;
        RECT 2131.450 2595.060 2144.150 2595.340 ;
        RECT 2132.850 2594.780 2142.750 2595.060 ;
        RECT 2133.940 2594.500 2141.660 2594.780 ;
        RECT 2134.790 2594.220 2140.810 2594.500 ;
        RECT 2135.300 2569.720 2140.300 2594.220 ;
        RECT 2028.365 2564.720 2140.300 2569.720 ;
        RECT 2028.365 2274.920 2033.365 2564.720 ;
        RECT 2028.315 2269.920 2033.415 2274.920 ;
      LAYER Metal3 ;
        RECT 2028.365 2274.920 2033.365 2274.965 ;
        RECT 2028.320 2269.920 2033.410 2274.920 ;
        RECT 2028.365 2269.875 2033.365 2269.920 ;
      LAYER Metal4 ;
        RECT 2028.365 2274.920 2033.365 2274.965 ;
        RECT 2028.320 2269.920 2033.410 2274.920 ;
        RECT 2028.365 2269.875 2033.365 2269.920 ;
      LAYER Metal5 ;
        RECT 2028.365 2274.920 2033.365 2274.965 ;
        RECT 1985.365 2269.920 2053.365 2274.920 ;
        RECT 2028.365 2269.875 2033.365 2269.920 ;
    END
  END vss_pad_n_4
  PIN vddcore0_pad_n_5
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal2 ;
        RECT 2001.660 2605.300 2011.160 2606.300 ;
        RECT 2014.060 2605.300 2024.310 2606.300 ;
        RECT 2025.910 2605.300 2036.160 2606.300 ;
        RECT 2039.440 2605.300 2049.690 2606.300 ;
        RECT 2051.290 2605.300 2061.540 2606.300 ;
        RECT 2064.440 2605.300 2073.940 2606.300 ;
        RECT 2001.660 2597.020 2073.940 2605.300 ;
        RECT 2009.610 2596.740 2065.990 2597.020 ;
        RECT 2015.810 2596.460 2059.790 2596.740 ;
        RECT 2020.650 2596.180 2054.950 2596.460 ;
        RECT 2024.420 2595.900 2051.180 2596.180 ;
        RECT 2027.370 2595.620 2048.230 2595.900 ;
        RECT 2029.660 2595.340 2045.940 2595.620 ;
        RECT 2031.450 2595.060 2044.150 2595.340 ;
        RECT 2032.850 2594.780 2042.750 2595.060 ;
        RECT 2033.940 2594.500 2041.660 2594.780 ;
        RECT 2034.790 2594.220 2040.810 2594.500 ;
        RECT 2035.300 2584.720 2040.300 2594.220 ;
        RECT 2005.365 2579.720 2040.300 2584.720 ;
        RECT 2005.365 2267.920 2010.365 2579.720 ;
        RECT 2005.315 2262.920 2010.415 2267.920 ;
      LAYER Metal3 ;
        RECT 2005.365 2267.920 2010.365 2267.965 ;
        RECT 2005.320 2262.920 2010.410 2267.920 ;
        RECT 2005.365 2262.875 2010.365 2262.920 ;
      LAYER Metal4 ;
        RECT 2005.365 2267.920 2010.365 2267.965 ;
        RECT 2005.320 2262.920 2010.410 2267.920 ;
        RECT 2005.365 2262.875 2010.365 2262.920 ;
      LAYER Metal5 ;
        RECT 2005.365 2267.920 2010.365 2267.965 ;
        RECT 1985.365 2262.920 2053.365 2267.920 ;
        RECT 2005.365 2262.875 2010.365 2262.920 ;
    END
  END vddcore0_pad_n_5
  PIN vss_pad_n_16
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal2 ;
        RECT 901.660 2605.300 911.160 2606.300 ;
        RECT 914.060 2605.300 924.310 2606.300 ;
        RECT 925.910 2605.300 936.160 2606.300 ;
        RECT 939.440 2605.300 949.690 2606.300 ;
        RECT 951.290 2605.300 961.540 2606.300 ;
        RECT 964.440 2605.300 973.940 2606.300 ;
        RECT 901.660 2597.020 973.940 2605.300 ;
        RECT 909.610 2596.740 965.990 2597.020 ;
        RECT 915.810 2596.460 959.790 2596.740 ;
        RECT 920.650 2596.180 954.950 2596.460 ;
        RECT 924.420 2595.900 951.180 2596.180 ;
        RECT 927.370 2595.620 948.230 2595.900 ;
        RECT 929.660 2595.340 945.940 2595.620 ;
        RECT 931.450 2595.060 944.150 2595.340 ;
        RECT 932.850 2594.780 942.750 2595.060 ;
        RECT 933.940 2594.500 941.660 2594.780 ;
        RECT 934.790 2594.220 940.810 2594.500 ;
        RECT 935.300 2274.920 940.300 2594.220 ;
        RECT 935.250 2269.920 940.350 2274.920 ;
      LAYER Metal3 ;
        RECT 935.300 2274.920 940.300 2274.965 ;
        RECT 935.255 2269.920 940.345 2274.920 ;
        RECT 935.300 2269.875 940.300 2269.920 ;
      LAYER Metal4 ;
        RECT 935.300 2274.920 940.300 2274.965 ;
        RECT 935.255 2269.920 940.345 2274.920 ;
        RECT 935.300 2269.875 940.300 2269.920 ;
      LAYER Metal5 ;
        RECT 935.300 2274.920 940.300 2274.965 ;
        RECT 915.300 2269.920 960.300 2274.920 ;
        RECT 935.300 2269.875 940.300 2269.920 ;
    END
  END vss_pad_n_16
  PIN vss_pad_n_18
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal2 ;
        RECT 701.660 2605.300 711.160 2606.300 ;
        RECT 714.060 2605.300 724.310 2606.300 ;
        RECT 725.910 2605.300 736.160 2606.300 ;
        RECT 739.440 2605.300 749.690 2606.300 ;
        RECT 751.290 2605.300 761.540 2606.300 ;
        RECT 764.440 2605.300 773.940 2606.300 ;
        RECT 701.660 2597.020 773.940 2605.300 ;
        RECT 709.610 2596.740 765.990 2597.020 ;
        RECT 715.810 2596.460 759.790 2596.740 ;
        RECT 720.650 2596.180 754.950 2596.460 ;
        RECT 724.420 2595.900 751.180 2596.180 ;
        RECT 727.370 2595.620 748.230 2595.900 ;
        RECT 729.660 2595.340 745.940 2595.620 ;
        RECT 731.450 2595.060 744.150 2595.340 ;
        RECT 732.850 2594.780 742.750 2595.060 ;
        RECT 733.940 2594.500 741.660 2594.780 ;
        RECT 734.790 2594.220 740.810 2594.500 ;
        RECT 735.450 2593.940 740.150 2594.220 ;
        RECT 735.970 2593.660 739.630 2593.940 ;
        RECT 736.200 2575.420 739.400 2593.660 ;
        RECT 736.150 2573.820 739.400 2575.420 ;
        RECT 737.800 2552.660 739.400 2573.820 ;
        RECT 737.750 2551.060 739.450 2552.660 ;
      LAYER Metal3 ;
        RECT 736.200 2575.420 737.800 2575.470 ;
        RECT 612.800 2573.820 737.800 2575.420 ;
        RECT 612.800 2280.540 614.400 2573.820 ;
        RECT 736.200 2573.770 737.800 2573.820 ;
        RECT 737.800 2552.660 739.400 2552.705 ;
        RECT 737.755 2551.060 739.445 2552.660 ;
        RECT 737.800 2551.015 739.400 2551.060 ;
        RECT 612.750 2278.940 614.450 2280.540 ;
      LAYER Metal4 ;
        RECT 737.800 2552.660 739.400 2552.705 ;
        RECT 737.755 2551.060 739.445 2552.660 ;
        RECT 737.800 2551.015 739.400 2551.060 ;
        RECT 612.800 2280.540 614.400 2280.585 ;
        RECT 612.755 2278.940 614.445 2280.540 ;
        RECT 612.800 2278.895 614.400 2278.940 ;
      LAYER Metal5 ;
        RECT 737.800 2552.660 739.400 2552.705 ;
        RECT 721.400 2551.060 745.800 2552.660 ;
        RECT 737.800 2551.015 739.400 2551.060 ;
        RECT 612.800 2280.540 614.400 2280.585 ;
        RECT 596.400 2278.940 620.800 2280.540 ;
        RECT 612.800 2278.895 614.400 2278.940 ;
    END
  END vss_pad_n_18
  PIN vddcore1_pad_n_19
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal2 ;
        RECT 601.660 2605.300 611.160 2606.300 ;
        RECT 614.060 2605.300 624.310 2606.300 ;
        RECT 625.910 2605.300 636.160 2606.300 ;
        RECT 639.440 2605.300 649.690 2606.300 ;
        RECT 651.290 2605.300 661.540 2606.300 ;
        RECT 664.440 2605.300 673.940 2606.300 ;
        RECT 601.660 2597.020 673.940 2605.300 ;
        RECT 609.610 2596.740 665.990 2597.020 ;
        RECT 615.810 2596.460 659.790 2596.740 ;
        RECT 620.650 2596.180 654.950 2596.460 ;
        RECT 624.420 2595.900 651.180 2596.180 ;
        RECT 627.370 2595.620 648.230 2595.900 ;
        RECT 629.660 2595.340 645.940 2595.620 ;
        RECT 631.450 2595.060 644.150 2595.340 ;
        RECT 632.850 2594.780 642.750 2595.060 ;
        RECT 633.940 2594.500 641.660 2594.780 ;
        RECT 634.790 2594.220 640.810 2594.500 ;
        RECT 635.450 2593.940 640.150 2594.220 ;
        RECT 635.970 2593.660 639.630 2593.940 ;
        RECT 636.200 2586.420 639.400 2593.660 ;
        RECT 636.150 2584.820 729.400 2586.420 ;
        RECT 727.800 2549.360 729.400 2584.820 ;
        RECT 727.750 2547.760 729.450 2549.360 ;
      LAYER Metal3 ;
        RECT 636.200 2586.420 637.800 2586.470 ;
        RECT 602.800 2584.820 637.800 2586.420 ;
        RECT 602.800 2277.240 604.400 2584.820 ;
        RECT 636.200 2584.770 637.800 2584.820 ;
        RECT 727.800 2549.360 729.400 2549.405 ;
        RECT 727.755 2547.760 729.445 2549.360 ;
        RECT 727.800 2547.715 729.400 2547.760 ;
        RECT 602.750 2275.640 604.450 2277.240 ;
      LAYER Metal4 ;
        RECT 727.800 2549.360 729.400 2549.405 ;
        RECT 727.755 2547.760 729.445 2549.360 ;
        RECT 727.800 2547.715 729.400 2547.760 ;
        RECT 602.800 2277.240 604.400 2277.285 ;
        RECT 602.755 2275.640 604.445 2277.240 ;
        RECT 602.800 2275.595 604.400 2275.640 ;
      LAYER Metal5 ;
        RECT 727.800 2549.360 729.400 2549.405 ;
        RECT 721.400 2547.760 745.800 2549.360 ;
        RECT 727.800 2547.715 729.400 2547.760 ;
        RECT 602.800 2277.240 604.400 2277.285 ;
        RECT 596.400 2275.640 620.800 2277.240 ;
        RECT 602.800 2275.595 604.400 2275.640 ;
    END
  END vddcore1_pad_n_19
  PIN vss_pad_w_2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal2 ;
        RECT 369.300 2365.990 378.580 2373.940 ;
        RECT 369.300 2364.440 378.860 2365.990 ;
        RECT 370.300 2361.540 378.860 2364.440 ;
        RECT 369.300 2359.790 378.860 2361.540 ;
        RECT 369.300 2354.950 379.140 2359.790 ;
        RECT 692.220 2358.600 693.820 2358.650 ;
        RECT 389.180 2357.000 693.820 2358.600 ;
        RECT 369.300 2351.290 379.420 2354.950 ;
        RECT 370.300 2351.180 379.420 2351.290 ;
        RECT 370.300 2349.690 379.700 2351.180 ;
        RECT 369.300 2348.230 379.700 2349.690 ;
        RECT 369.300 2345.940 379.980 2348.230 ;
        RECT 369.300 2344.150 380.260 2345.940 ;
        RECT 369.300 2342.750 380.540 2344.150 ;
        RECT 369.300 2341.660 380.820 2342.750 ;
        RECT 369.300 2340.810 381.100 2341.660 ;
        RECT 369.300 2340.150 381.380 2340.810 ;
        RECT 369.300 2339.630 381.660 2340.150 ;
        RECT 369.300 2339.440 381.940 2339.630 ;
        RECT 370.300 2339.400 381.940 2339.440 ;
        RECT 389.180 2339.400 390.780 2357.000 ;
        RECT 692.220 2356.950 693.820 2357.000 ;
        RECT 370.300 2336.200 390.780 2339.400 ;
        RECT 370.300 2336.160 381.940 2336.200 ;
        RECT 369.300 2335.970 381.940 2336.160 ;
        RECT 369.300 2335.450 381.660 2335.970 ;
        RECT 369.300 2334.790 381.380 2335.450 ;
        RECT 369.300 2333.940 381.100 2334.790 ;
        RECT 369.300 2332.850 380.820 2333.940 ;
        RECT 369.300 2331.450 380.540 2332.850 ;
        RECT 369.300 2329.660 380.260 2331.450 ;
        RECT 369.300 2327.370 379.980 2329.660 ;
        RECT 369.300 2325.910 379.700 2327.370 ;
        RECT 370.300 2324.420 379.700 2325.910 ;
        RECT 370.300 2324.310 379.420 2324.420 ;
        RECT 369.300 2320.650 379.420 2324.310 ;
        RECT 369.300 2315.810 379.140 2320.650 ;
        RECT 369.300 2314.060 378.860 2315.810 ;
        RECT 370.300 2311.160 378.860 2314.060 ;
        RECT 369.300 2309.610 378.860 2311.160 ;
        RECT 369.300 2301.660 378.580 2309.610 ;
        RECT 389.180 2253.600 390.780 2336.200 ;
        RECT 421.220 2253.600 422.820 2253.650 ;
        RECT 389.180 2252.000 422.820 2253.600 ;
        RECT 421.220 2251.950 422.820 2252.000 ;
      LAYER Metal3 ;
        RECT 692.220 2358.600 693.820 2358.645 ;
        RECT 692.175 2357.000 693.865 2358.600 ;
        RECT 692.220 2356.955 693.820 2357.000 ;
        RECT 421.220 2253.600 422.820 2253.645 ;
        RECT 421.175 2252.000 422.865 2253.600 ;
        RECT 421.220 2251.955 422.820 2252.000 ;
      LAYER Metal4 ;
        RECT 692.220 2358.600 693.820 2365.000 ;
        RECT 692.175 2357.000 693.865 2358.600 ;
        RECT 692.220 2350.600 693.820 2357.000 ;
        RECT 421.220 2253.600 422.820 2260.000 ;
        RECT 421.175 2252.000 422.865 2253.600 ;
        RECT 421.220 2245.600 422.820 2252.000 ;
    END
  END vss_pad_w_2
  PIN vss_pad_w_4
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal2 ;
        RECT 369.300 2165.990 378.580 2173.940 ;
        RECT 369.300 2164.440 378.860 2165.990 ;
        RECT 370.300 2161.540 378.860 2164.440 ;
        RECT 369.300 2159.790 378.860 2161.540 ;
        RECT 369.300 2154.950 379.140 2159.790 ;
        RECT 369.300 2151.290 379.420 2154.950 ;
        RECT 370.300 2151.180 379.420 2151.290 ;
        RECT 370.300 2149.690 379.700 2151.180 ;
        RECT 369.300 2148.230 379.700 2149.690 ;
        RECT 369.300 2145.940 379.980 2148.230 ;
        RECT 369.300 2144.150 380.260 2145.940 ;
        RECT 369.300 2142.750 380.540 2144.150 ;
        RECT 369.300 2141.660 380.820 2142.750 ;
        RECT 369.300 2140.810 381.100 2141.660 ;
        RECT 369.300 2140.300 381.380 2140.810 ;
        RECT 369.300 2139.440 410.880 2140.300 ;
        RECT 370.300 2136.160 410.880 2139.440 ;
        RECT 369.300 2135.300 410.880 2136.160 ;
        RECT 369.300 2134.790 381.380 2135.300 ;
        RECT 369.300 2133.940 381.100 2134.790 ;
        RECT 369.300 2132.850 380.820 2133.940 ;
        RECT 369.300 2131.450 380.540 2132.850 ;
        RECT 369.300 2129.660 380.260 2131.450 ;
        RECT 369.300 2127.370 379.980 2129.660 ;
        RECT 369.300 2125.910 379.700 2127.370 ;
        RECT 370.300 2124.420 379.700 2125.910 ;
        RECT 370.300 2124.310 379.420 2124.420 ;
        RECT 369.300 2120.650 379.420 2124.310 ;
        RECT 369.300 2115.810 379.140 2120.650 ;
        RECT 369.300 2114.060 378.860 2115.810 ;
        RECT 370.300 2111.160 378.860 2114.060 ;
        RECT 369.300 2109.610 378.860 2111.160 ;
        RECT 369.300 2101.660 378.580 2109.610 ;
        RECT 405.880 2033.365 410.880 2135.300 ;
        RECT 698.200 2033.365 703.200 2033.415 ;
        RECT 405.880 2028.365 703.200 2033.365 ;
        RECT 698.200 2028.315 703.200 2028.365 ;
      LAYER Metal3 ;
        RECT 698.200 2033.365 703.200 2033.410 ;
        RECT 698.155 2028.365 703.245 2033.365 ;
        RECT 698.200 2028.320 703.200 2028.365 ;
      LAYER Metal4 ;
        RECT 698.200 2033.365 703.200 2053.365 ;
        RECT 698.155 2028.365 703.245 2033.365 ;
        RECT 698.200 1988.365 703.200 2028.365 ;
    END
  END vss_pad_w_4
  PIN vddcore0_pad_w_5
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal2 ;
        RECT 369.300 2065.990 378.580 2073.940 ;
        RECT 369.300 2064.440 378.860 2065.990 ;
        RECT 370.300 2061.540 378.860 2064.440 ;
        RECT 369.300 2059.790 378.860 2061.540 ;
        RECT 369.300 2054.950 379.140 2059.790 ;
        RECT 369.300 2051.290 379.420 2054.950 ;
        RECT 370.300 2051.180 379.420 2051.290 ;
        RECT 370.300 2049.690 379.700 2051.180 ;
        RECT 369.300 2048.230 379.700 2049.690 ;
        RECT 369.300 2045.940 379.980 2048.230 ;
        RECT 369.300 2044.150 380.260 2045.940 ;
        RECT 369.300 2042.750 380.540 2044.150 ;
        RECT 369.300 2041.660 380.820 2042.750 ;
        RECT 369.300 2040.810 381.100 2041.660 ;
        RECT 369.300 2040.300 381.380 2040.810 ;
        RECT 369.300 2039.440 395.880 2040.300 ;
        RECT 370.300 2036.160 395.880 2039.440 ;
        RECT 369.300 2035.300 395.880 2036.160 ;
        RECT 369.300 2034.790 381.380 2035.300 ;
        RECT 369.300 2033.940 381.100 2034.790 ;
        RECT 369.300 2032.850 380.820 2033.940 ;
        RECT 369.300 2031.450 380.540 2032.850 ;
        RECT 369.300 2029.660 380.260 2031.450 ;
        RECT 369.300 2027.370 379.980 2029.660 ;
        RECT 369.300 2025.910 379.700 2027.370 ;
        RECT 370.300 2024.420 379.700 2025.910 ;
        RECT 370.300 2024.310 379.420 2024.420 ;
        RECT 369.300 2020.650 379.420 2024.310 ;
        RECT 369.300 2015.810 379.140 2020.650 ;
        RECT 369.300 2014.060 378.860 2015.810 ;
        RECT 370.300 2011.160 378.860 2014.060 ;
        RECT 369.300 2009.610 378.860 2011.160 ;
        RECT 390.880 2013.365 395.880 2035.300 ;
        RECT 705.200 2013.365 710.200 2013.415 ;
        RECT 369.300 2001.660 378.580 2009.610 ;
        RECT 390.880 2008.365 710.200 2013.365 ;
        RECT 705.200 2008.315 710.200 2008.365 ;
      LAYER Metal3 ;
        RECT 705.200 2013.365 710.200 2013.410 ;
        RECT 705.155 2008.365 710.245 2013.365 ;
        RECT 705.200 2008.320 710.200 2008.365 ;
      LAYER Metal4 ;
        RECT 705.200 2013.365 710.200 2053.365 ;
        RECT 705.155 2008.365 710.245 2013.365 ;
        RECT 705.200 1988.365 710.200 2008.365 ;
    END
  END vddcore0_pad_w_5
  PIN vss_pad_w_16
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal2 ;
        RECT 369.300 965.990 378.580 973.940 ;
        RECT 369.300 964.440 378.860 965.990 ;
        RECT 370.300 961.540 378.860 964.440 ;
        RECT 369.300 959.790 378.860 961.540 ;
        RECT 369.300 954.950 379.140 959.790 ;
        RECT 369.300 951.290 379.420 954.950 ;
        RECT 370.300 951.180 379.420 951.290 ;
        RECT 370.300 949.690 379.700 951.180 ;
        RECT 369.300 948.230 379.700 949.690 ;
        RECT 369.300 945.940 379.980 948.230 ;
        RECT 369.300 944.150 380.260 945.940 ;
        RECT 369.300 942.750 380.540 944.150 ;
        RECT 369.300 941.660 380.820 942.750 ;
        RECT 369.300 940.810 381.100 941.660 ;
        RECT 369.300 940.300 381.380 940.810 ;
        RECT 698.200 940.300 703.200 940.350 ;
        RECT 369.300 939.440 703.200 940.300 ;
        RECT 370.300 936.160 703.200 939.440 ;
        RECT 369.300 935.300 703.200 936.160 ;
        RECT 369.300 934.790 381.380 935.300 ;
        RECT 698.200 935.250 703.200 935.300 ;
        RECT 369.300 933.940 381.100 934.790 ;
        RECT 369.300 932.850 380.820 933.940 ;
        RECT 369.300 931.450 380.540 932.850 ;
        RECT 369.300 929.660 380.260 931.450 ;
        RECT 369.300 927.370 379.980 929.660 ;
        RECT 369.300 925.910 379.700 927.370 ;
        RECT 370.300 924.420 379.700 925.910 ;
        RECT 370.300 924.310 379.420 924.420 ;
        RECT 369.300 920.650 379.420 924.310 ;
        RECT 369.300 915.810 379.140 920.650 ;
        RECT 369.300 914.060 378.860 915.810 ;
        RECT 370.300 911.160 378.860 914.060 ;
        RECT 369.300 909.610 378.860 911.160 ;
        RECT 369.300 901.660 378.580 909.610 ;
      LAYER Metal3 ;
        RECT 698.200 940.300 703.200 940.345 ;
        RECT 698.155 935.300 703.245 940.300 ;
        RECT 698.200 935.255 703.200 935.300 ;
      LAYER Metal4 ;
        RECT 698.200 940.300 703.200 960.300 ;
        RECT 698.155 935.300 703.245 940.300 ;
        RECT 698.200 915.300 703.200 935.300 ;
    END
  END vss_pad_w_16
  PIN vss_pad_w_18
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal2 ;
        RECT 369.300 765.990 378.580 773.940 ;
        RECT 369.300 764.440 378.860 765.990 ;
        RECT 370.300 761.540 378.860 764.440 ;
        RECT 369.300 759.790 378.860 761.540 ;
        RECT 369.300 754.950 379.140 759.790 ;
        RECT 369.300 751.290 379.420 754.950 ;
        RECT 370.300 751.180 379.420 751.290 ;
        RECT 370.300 749.690 379.700 751.180 ;
        RECT 369.300 748.230 379.700 749.690 ;
        RECT 369.300 745.940 379.980 748.230 ;
        RECT 369.300 744.150 380.260 745.940 ;
        RECT 369.300 742.750 380.540 744.150 ;
        RECT 369.300 741.660 380.820 742.750 ;
        RECT 369.300 740.810 381.100 741.660 ;
        RECT 369.300 740.150 381.380 740.810 ;
        RECT 369.300 739.630 381.660 740.150 ;
        RECT 369.300 739.440 381.940 739.630 ;
        RECT 370.300 739.400 381.940 739.440 ;
        RECT 370.300 737.800 412.780 739.400 ;
        RECT 421.220 737.800 422.820 737.850 ;
        RECT 370.300 736.200 401.780 737.800 ;
        RECT 411.180 736.200 422.820 737.800 ;
        RECT 370.300 736.160 381.940 736.200 ;
        RECT 369.300 735.970 381.940 736.160 ;
        RECT 400.180 736.150 401.780 736.200 ;
        RECT 421.220 736.150 422.820 736.200 ;
        RECT 369.300 735.450 381.660 735.970 ;
        RECT 369.300 734.790 381.380 735.450 ;
        RECT 369.300 733.940 381.100 734.790 ;
        RECT 369.300 732.850 380.820 733.940 ;
        RECT 369.300 731.450 380.540 732.850 ;
        RECT 369.300 729.660 380.260 731.450 ;
        RECT 369.300 727.370 379.980 729.660 ;
        RECT 369.300 725.910 379.700 727.370 ;
        RECT 370.300 724.420 379.700 725.910 ;
        RECT 370.300 724.310 379.420 724.420 ;
        RECT 369.300 720.650 379.420 724.310 ;
        RECT 369.300 715.810 379.140 720.650 ;
        RECT 369.300 714.060 378.860 715.810 ;
        RECT 370.300 711.160 378.860 714.060 ;
        RECT 369.300 709.610 378.860 711.160 ;
        RECT 369.300 701.660 378.580 709.610 ;
      LAYER Metal3 ;
        RECT 421.220 737.800 422.820 737.845 ;
        RECT 400.130 736.200 401.830 737.800 ;
        RECT 421.175 736.200 422.865 737.800 ;
        RECT 400.180 614.400 401.780 736.200 ;
        RECT 421.220 736.155 422.820 736.200 ;
        RECT 692.220 614.400 693.820 614.450 ;
        RECT 400.180 612.800 693.820 614.400 ;
        RECT 692.220 612.750 693.820 612.800 ;
      LAYER Metal4 ;
        RECT 421.220 737.800 422.820 744.200 ;
        RECT 421.175 736.200 422.865 737.800 ;
        RECT 421.220 721.400 422.820 736.200 ;
        RECT 692.220 614.400 693.820 620.800 ;
        RECT 692.175 612.800 693.865 614.400 ;
        RECT 692.220 596.400 693.820 612.800 ;
    END
  END vss_pad_w_18
  PIN vddcore2_pad_w_19
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal2 ;
        RECT 424.520 729.400 426.120 729.450 ;
        RECT 389.180 727.800 426.120 729.400 ;
        RECT 369.300 665.990 378.580 673.940 ;
        RECT 369.300 664.440 378.860 665.990 ;
        RECT 370.300 661.540 378.860 664.440 ;
        RECT 369.300 659.790 378.860 661.540 ;
        RECT 369.300 654.950 379.140 659.790 ;
        RECT 369.300 651.290 379.420 654.950 ;
        RECT 370.300 651.180 379.420 651.290 ;
        RECT 370.300 649.690 379.700 651.180 ;
        RECT 369.300 648.230 379.700 649.690 ;
        RECT 369.300 645.940 379.980 648.230 ;
        RECT 369.300 644.150 380.260 645.940 ;
        RECT 369.300 642.750 380.540 644.150 ;
        RECT 369.300 641.660 380.820 642.750 ;
        RECT 369.300 640.810 381.100 641.660 ;
        RECT 369.300 640.150 381.380 640.810 ;
        RECT 369.300 639.630 381.660 640.150 ;
        RECT 369.300 639.440 381.940 639.630 ;
        RECT 370.300 639.400 381.940 639.440 ;
        RECT 389.180 639.400 390.780 727.800 ;
        RECT 424.520 727.750 426.120 727.800 ;
        RECT 370.300 636.200 390.780 639.400 ;
        RECT 370.300 636.160 381.940 636.200 ;
        RECT 369.300 635.970 381.940 636.160 ;
        RECT 389.180 636.150 390.780 636.200 ;
        RECT 369.300 635.450 381.660 635.970 ;
        RECT 369.300 634.790 381.380 635.450 ;
        RECT 369.300 633.940 381.100 634.790 ;
        RECT 369.300 632.850 380.820 633.940 ;
        RECT 369.300 631.450 380.540 632.850 ;
        RECT 369.300 629.660 380.260 631.450 ;
        RECT 369.300 627.370 379.980 629.660 ;
        RECT 369.300 625.910 379.700 627.370 ;
        RECT 370.300 624.420 379.700 625.910 ;
        RECT 370.300 624.310 379.420 624.420 ;
        RECT 369.300 620.650 379.420 624.310 ;
        RECT 369.300 615.810 379.140 620.650 ;
        RECT 369.300 614.060 378.860 615.810 ;
        RECT 370.300 611.160 378.860 614.060 ;
        RECT 369.300 609.610 378.860 611.160 ;
        RECT 369.300 601.660 378.580 609.610 ;
      LAYER Metal3 ;
        RECT 424.520 729.400 426.120 729.445 ;
        RECT 424.475 727.800 426.165 729.400 ;
        RECT 424.520 727.755 426.120 727.800 ;
        RECT 389.130 636.200 390.830 637.800 ;
        RECT 389.180 604.400 390.780 636.200 ;
        RECT 695.520 604.400 697.120 604.450 ;
        RECT 389.180 602.800 697.120 604.400 ;
        RECT 695.520 602.750 697.120 602.800 ;
      LAYER Metal4 ;
        RECT 424.520 729.400 426.120 744.200 ;
        RECT 424.475 727.800 426.165 729.400 ;
        RECT 424.520 721.400 426.120 727.800 ;
        RECT 695.520 604.400 697.120 620.800 ;
        RECT 695.475 602.800 697.165 604.400 ;
        RECT 695.520 596.400 697.120 602.800 ;
    END
  END vddcore2_pad_w_19
  PIN loop_pad_s_6
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1037.610 383.900 1037.990 388.680 ;
        RECT 1037.600 383.620 1038.000 383.900 ;
        RECT 1037.550 383.340 1038.050 383.620 ;
        RECT 1037.480 383.060 1038.120 383.340 ;
        RECT 1037.380 382.780 1038.220 383.060 ;
        RECT 1037.270 382.500 1038.330 382.780 ;
        RECT 1037.120 382.220 1038.480 382.500 ;
        RECT 1036.920 381.940 1038.680 382.220 ;
        RECT 1036.680 381.660 1038.920 381.940 ;
        RECT 1036.360 381.380 1039.240 381.660 ;
        RECT 1035.950 381.100 1039.650 381.380 ;
        RECT 1035.430 380.820 1040.170 381.100 ;
        RECT 1034.760 380.540 1040.840 380.820 ;
        RECT 1033.910 380.260 1041.690 380.540 ;
        RECT 1032.810 379.980 1042.790 380.260 ;
        RECT 1031.400 379.700 1044.200 379.980 ;
        RECT 1029.600 379.420 1046.000 379.700 ;
        RECT 1027.280 379.140 1048.320 379.420 ;
        RECT 1024.320 378.860 1051.280 379.140 ;
        RECT 1020.520 378.580 1055.080 378.860 ;
        RECT 1015.640 370.300 1059.960 378.580 ;
        RECT 1015.640 369.300 1018.180 370.300 ;
        RECT 1021.320 369.300 1023.860 370.300 ;
        RECT 1027.000 369.300 1029.540 370.300 ;
        RECT 1032.680 369.300 1035.220 370.300 ;
        RECT 1040.380 369.300 1042.920 370.300 ;
        RECT 1046.060 369.300 1048.600 370.300 ;
        RECT 1051.740 369.300 1054.280 370.300 ;
        RECT 1057.420 369.300 1059.960 370.300 ;
    END
  END loop_pad_s_6
  PIN loop_pad_s_7
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1137.610 383.900 1137.990 388.680 ;
        RECT 1137.600 383.620 1138.000 383.900 ;
        RECT 1137.550 383.340 1138.050 383.620 ;
        RECT 1137.480 383.060 1138.120 383.340 ;
        RECT 1137.380 382.780 1138.220 383.060 ;
        RECT 1137.270 382.500 1138.330 382.780 ;
        RECT 1137.120 382.220 1138.480 382.500 ;
        RECT 1136.920 381.940 1138.680 382.220 ;
        RECT 1136.680 381.660 1138.920 381.940 ;
        RECT 1136.360 381.380 1139.240 381.660 ;
        RECT 1135.950 381.100 1139.650 381.380 ;
        RECT 1135.430 380.820 1140.170 381.100 ;
        RECT 1134.760 380.540 1140.840 380.820 ;
        RECT 1133.910 380.260 1141.690 380.540 ;
        RECT 1132.810 379.980 1142.790 380.260 ;
        RECT 1131.400 379.700 1144.200 379.980 ;
        RECT 1129.600 379.420 1146.000 379.700 ;
        RECT 1127.280 379.140 1148.320 379.420 ;
        RECT 1124.320 378.860 1151.280 379.140 ;
        RECT 1120.520 378.580 1155.080 378.860 ;
        RECT 1115.640 370.300 1159.960 378.580 ;
        RECT 1115.640 369.300 1118.180 370.300 ;
        RECT 1121.320 369.300 1123.860 370.300 ;
        RECT 1127.000 369.300 1129.540 370.300 ;
        RECT 1132.680 369.300 1135.220 370.300 ;
        RECT 1140.380 369.300 1142.920 370.300 ;
        RECT 1146.060 369.300 1148.600 370.300 ;
        RECT 1151.740 369.300 1154.280 370.300 ;
        RECT 1157.420 369.300 1159.960 370.300 ;
    END
  END loop_pad_s_7
  PIN tie_pad_n_12
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1315.640 2605.300 1318.180 2606.300 ;
        RECT 1321.320 2605.300 1323.860 2606.300 ;
        RECT 1327.000 2605.300 1329.540 2606.300 ;
        RECT 1332.680 2605.300 1335.220 2606.300 ;
        RECT 1340.380 2605.300 1342.920 2606.300 ;
        RECT 1346.060 2605.300 1348.600 2606.300 ;
        RECT 1351.740 2605.300 1354.280 2606.300 ;
        RECT 1357.420 2605.300 1359.960 2606.300 ;
        RECT 1315.640 2597.020 1359.960 2605.300 ;
        RECT 1320.520 2596.740 1355.080 2597.020 ;
        RECT 1324.320 2596.460 1351.280 2596.740 ;
        RECT 1327.280 2596.180 1348.320 2596.460 ;
        RECT 1329.600 2595.900 1346.000 2596.180 ;
        RECT 1331.400 2595.620 1344.200 2595.900 ;
        RECT 1332.810 2595.340 1342.790 2595.620 ;
        RECT 1333.910 2595.060 1341.690 2595.340 ;
        RECT 1334.760 2594.780 1340.840 2595.060 ;
        RECT 1335.430 2594.500 1340.170 2594.780 ;
        RECT 1335.950 2594.220 1339.650 2594.500 ;
        RECT 1336.360 2593.940 1339.240 2594.220 ;
        RECT 1336.680 2593.660 1338.920 2593.940 ;
        RECT 1336.920 2593.380 1338.680 2593.660 ;
        RECT 1337.120 2593.100 1338.480 2593.380 ;
        RECT 1337.270 2592.820 1338.330 2593.100 ;
        RECT 1337.380 2592.540 1338.220 2592.820 ;
        RECT 1337.480 2592.260 1338.120 2592.540 ;
        RECT 1337.550 2591.980 1338.050 2592.260 ;
        RECT 1337.600 2591.700 1338.000 2591.980 ;
        RECT 1337.610 2589.300 1337.990 2591.700 ;
        RECT 1411.685 2589.300 1412.065 2605.300 ;
        RECT 1337.610 2588.920 1412.065 2589.300 ;
    END
  END tie_pad_n_12
  PIN ta_pad_n_13
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1215.640 2605.300 1218.180 2606.300 ;
        RECT 1221.320 2605.300 1223.860 2606.300 ;
        RECT 1227.000 2605.300 1229.540 2606.300 ;
        RECT 1232.680 2605.300 1235.220 2606.300 ;
        RECT 1240.380 2605.300 1242.920 2606.300 ;
        RECT 1246.060 2605.300 1248.600 2606.300 ;
        RECT 1251.740 2605.300 1254.280 2606.300 ;
        RECT 1257.420 2605.300 1259.960 2606.300 ;
        RECT 1215.640 2597.020 1259.960 2605.300 ;
        RECT 1220.520 2596.740 1255.080 2597.020 ;
        RECT 1224.320 2596.460 1251.280 2596.740 ;
        RECT 1227.280 2596.180 1248.320 2596.460 ;
        RECT 1229.600 2595.900 1246.000 2596.180 ;
        RECT 1231.400 2595.620 1244.200 2595.900 ;
        RECT 1232.810 2595.340 1242.790 2595.620 ;
        RECT 1233.910 2595.060 1241.690 2595.340 ;
        RECT 1234.760 2594.780 1240.840 2595.060 ;
        RECT 1235.430 2594.500 1240.170 2594.780 ;
        RECT 1235.950 2594.220 1239.650 2594.500 ;
        RECT 1236.360 2593.940 1239.240 2594.220 ;
        RECT 1236.680 2593.660 1238.920 2593.940 ;
        RECT 1236.920 2593.380 1238.680 2593.660 ;
        RECT 1237.120 2593.100 1238.480 2593.380 ;
        RECT 1237.270 2592.820 1238.330 2593.100 ;
        RECT 1237.380 2592.540 1238.220 2592.820 ;
        RECT 1237.480 2592.260 1238.120 2592.540 ;
        RECT 1237.550 2591.980 1238.050 2592.260 ;
        RECT 1237.600 2591.700 1238.000 2591.980 ;
        RECT 1237.610 2587.300 1237.990 2591.700 ;
        RECT 1469.700 2587.300 1470.080 2605.300 ;
        RECT 1237.610 2586.920 1470.080 2587.300 ;
    END
  END ta_pad_n_13
  PIN toe_pad_n_14
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1115.640 2605.300 1118.180 2606.300 ;
        RECT 1121.320 2605.300 1123.860 2606.300 ;
        RECT 1127.000 2605.300 1129.540 2606.300 ;
        RECT 1132.680 2605.300 1135.220 2606.300 ;
        RECT 1140.380 2605.300 1142.920 2606.300 ;
        RECT 1146.060 2605.300 1148.600 2606.300 ;
        RECT 1151.740 2605.300 1154.280 2606.300 ;
        RECT 1157.420 2605.300 1159.960 2606.300 ;
        RECT 1115.640 2597.020 1159.960 2605.300 ;
        RECT 1120.520 2596.740 1155.080 2597.020 ;
        RECT 1124.320 2596.460 1151.280 2596.740 ;
        RECT 1127.280 2596.180 1148.320 2596.460 ;
        RECT 1129.600 2595.900 1146.000 2596.180 ;
        RECT 1131.400 2595.620 1144.200 2595.900 ;
        RECT 1132.810 2595.340 1142.790 2595.620 ;
        RECT 1133.910 2595.060 1141.690 2595.340 ;
        RECT 1134.760 2594.780 1140.840 2595.060 ;
        RECT 1135.430 2594.500 1140.170 2594.780 ;
        RECT 1135.950 2594.220 1139.650 2594.500 ;
        RECT 1136.360 2593.940 1139.240 2594.220 ;
        RECT 1136.680 2593.660 1138.920 2593.940 ;
        RECT 1136.920 2593.380 1138.680 2593.660 ;
        RECT 1137.120 2593.100 1138.480 2593.380 ;
        RECT 1137.270 2592.820 1138.330 2593.100 ;
        RECT 1137.380 2592.540 1138.220 2592.820 ;
        RECT 1137.480 2592.260 1138.120 2592.540 ;
        RECT 1137.550 2591.980 1138.050 2592.260 ;
        RECT 1137.600 2591.700 1138.000 2591.980 ;
        RECT 1137.610 2585.300 1137.990 2591.700 ;
        RECT 1470.430 2585.300 1470.810 2605.300 ;
        RECT 1137.610 2584.920 1470.810 2585.300 ;
    END
  END toe_pad_n_14
  PIN ty_pad_n_15
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1015.640 2605.300 1018.180 2606.300 ;
        RECT 1021.320 2605.300 1023.860 2606.300 ;
        RECT 1027.000 2605.300 1029.540 2606.300 ;
        RECT 1032.680 2605.300 1035.220 2606.300 ;
        RECT 1040.380 2605.300 1042.920 2606.300 ;
        RECT 1046.060 2605.300 1048.600 2606.300 ;
        RECT 1051.740 2605.300 1054.280 2606.300 ;
        RECT 1057.420 2605.300 1059.960 2606.300 ;
        RECT 1015.640 2597.020 1059.960 2605.300 ;
        RECT 1020.520 2596.740 1055.080 2597.020 ;
        RECT 1024.320 2596.460 1051.280 2596.740 ;
        RECT 1027.280 2596.180 1048.320 2596.460 ;
        RECT 1029.600 2595.900 1046.000 2596.180 ;
        RECT 1031.400 2595.620 1044.200 2595.900 ;
        RECT 1032.810 2595.340 1042.790 2595.620 ;
        RECT 1033.910 2595.060 1041.690 2595.340 ;
        RECT 1034.760 2594.780 1040.840 2595.060 ;
        RECT 1035.430 2594.500 1040.170 2594.780 ;
        RECT 1035.950 2594.220 1039.650 2594.500 ;
        RECT 1036.360 2593.940 1039.240 2594.220 ;
        RECT 1036.680 2593.660 1038.920 2593.940 ;
        RECT 1036.920 2593.380 1038.680 2593.660 ;
        RECT 1037.120 2593.100 1038.480 2593.380 ;
        RECT 1037.270 2592.820 1038.330 2593.100 ;
        RECT 1037.380 2592.540 1038.220 2592.820 ;
        RECT 1037.480 2592.260 1038.120 2592.540 ;
        RECT 1037.550 2591.980 1038.050 2592.260 ;
        RECT 1037.600 2591.700 1038.000 2591.980 ;
        RECT 1037.610 2583.300 1037.990 2591.700 ;
        RECT 1471.160 2583.300 1471.540 2605.300 ;
        RECT 1037.610 2582.920 1471.540 2583.300 ;
    END
  END ty_pad_n_15
END wiring
END LIBRARY

