`default_nettype none

(* blackbox *)
module tt_logo (
    inout wire dummy
);

endmodule
