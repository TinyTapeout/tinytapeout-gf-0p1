`default_nettype none

(* blackbox *)
module loopback (
    inout wire A,
    inout wire B
);

endmodule
