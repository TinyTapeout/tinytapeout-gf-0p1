magic
tech gf180mcuD
magscale 1 10
timestamp 1757383304
<< metal2 >>
rect 127240 518884 127880 520332
rect 127230 518564 127240 518884
rect 127560 518564 144880 518884
rect 144560 509872 144880 518564
rect 147240 515884 147880 520332
rect 147230 515564 147240 515884
rect 147560 510532 147880 515884
rect 147550 510212 147560 510532
rect 147880 510212 147890 510532
rect 144550 509552 144560 509872
rect 144880 509552 144890 509872
rect 138444 471720 138764 471730
rect 76236 471400 138444 471720
rect 76236 467880 76556 471400
rect 138444 471390 138764 471400
rect 74788 467240 76556 467880
rect 76236 450720 76556 467240
rect 187060 454984 188060 520444
rect 207522 518260 207598 519940
rect 227522 518660 227598 519940
rect 247522 519060 247598 519940
rect 267522 519460 267598 519940
rect 282337 519460 282413 521060
rect 267522 519384 282413 519460
rect 293940 519060 294016 521060
rect 247522 518984 294016 519060
rect 294086 518660 294162 521060
rect 227522 518584 294162 518660
rect 294232 518260 294308 521060
rect 407060 518544 408060 520444
rect 207522 518184 294308 518260
rect 405673 517544 408060 518544
rect 187050 453984 187060 454984
rect 188060 453984 188070 454984
rect 405673 453584 406673 517544
rect 427060 515544 428060 520444
rect 467240 518884 467880 520332
rect 408673 514544 428060 515544
rect 450400 518564 471720 518884
rect 408673 454984 409673 514544
rect 450400 510532 450720 518564
rect 450390 510212 450400 510532
rect 450720 510212 450730 510532
rect 471400 456332 471720 518564
rect 518564 467880 518884 467890
rect 518884 467560 520332 467880
rect 518564 467240 520332 467560
rect 471390 456012 471400 456332
rect 471720 456012 471730 456332
rect 408663 453984 408673 454984
rect 409673 453984 409683 454984
rect 405663 452584 405673 453584
rect 406673 452584 406683 453584
rect 84244 450720 84564 450730
rect 76236 450400 84244 450720
rect 84244 450390 84564 450400
rect 510000 450560 510320 450570
rect 518564 450560 518884 467240
rect 510320 450240 518884 450560
rect 510000 450230 510320 450240
rect 515564 447880 515884 447890
rect 510660 447560 510980 447570
rect 515884 447560 520332 447880
rect 510980 447240 520332 447560
rect 510660 447230 510980 447240
rect 74676 427060 80576 428060
rect 79576 409673 80576 427060
rect 139640 409673 140640 409683
rect 79576 408673 139640 409673
rect 139640 408663 140640 408673
rect 454544 408060 455544 408070
rect 74676 407060 77576 408060
rect 76576 406673 77576 407060
rect 455544 407060 520444 408060
rect 454544 407050 455544 407060
rect 141040 406673 142040 406683
rect 76576 405673 141040 406673
rect 141040 405663 142040 405673
rect 453144 189447 454144 189457
rect 454144 188447 518544 189447
rect 453144 188437 454144 188447
rect 139640 188060 140640 188070
rect 74676 187060 139640 188060
rect 517544 188060 518544 188447
rect 517544 187060 520444 188060
rect 139640 187050 140640 187060
rect 454544 186447 455544 186457
rect 455544 185447 515544 186447
rect 454544 185437 455544 185447
rect 514544 168060 515544 185447
rect 514544 167060 520444 168060
rect 84244 147880 84564 147890
rect 74788 147560 84244 147880
rect 74788 147240 79236 147560
rect 84244 147550 84564 147560
rect 79236 147230 79556 147240
rect 84904 144880 85224 144890
rect 76236 144560 84904 144880
rect 76236 127880 76556 144560
rect 84904 144550 85224 144560
rect 510660 144720 510980 144730
rect 510980 144400 518884 144720
rect 510660 144390 510980 144400
rect 188437 141488 188447 142488
rect 189447 141488 189457 142488
rect 185437 140088 185447 141088
rect 186447 140088 186457 141088
rect 123390 138556 123400 138876
rect 123720 138556 123730 138876
rect 74788 127560 76556 127880
rect 74788 127240 76236 127560
rect 76236 127230 76556 127240
rect 123400 76556 123720 138556
rect 144390 84244 144400 84564
rect 144720 84244 144730 84564
rect 144400 76556 144720 84244
rect 185447 80576 186447 140088
rect 123400 76236 144720 76556
rect 167060 79576 186447 80576
rect 127240 74788 127880 76236
rect 167060 74676 168060 79576
rect 188447 77576 189447 141488
rect 407050 140088 407060 141088
rect 408060 140088 408070 141088
rect 187060 76576 189447 77576
rect 187060 74676 188060 76576
rect 207522 75180 207598 76136
rect 227522 75180 227598 76136
rect 407060 74676 408060 140088
rect 518564 127880 518884 144400
rect 518564 127240 520332 127880
rect 456460 123720 456780 123730
rect 518564 123720 518884 127240
rect 456780 123400 518884 123720
rect 456460 123390 456780 123400
rect 450230 85690 450240 86010
rect 450560 85690 450570 86010
rect 447230 85030 447240 85350
rect 447560 85030 447570 85350
rect 447240 79236 447560 85030
rect 447880 79236 447890 79556
rect 447240 74788 447880 79236
rect 450240 76556 450560 85690
rect 450240 76236 467560 76556
rect 467880 76236 467890 76556
rect 467240 74788 467880 76236
<< via2 >>
rect 127240 518564 127560 518884
rect 147240 515564 147560 515884
rect 147560 510212 147880 510532
rect 144560 509552 144880 509872
rect 138444 471400 138764 471720
rect 187060 453984 188060 454984
rect 450400 510212 450720 510532
rect 518564 467560 518884 467880
rect 471400 456012 471720 456332
rect 408673 453984 409673 454984
rect 405673 452584 406673 453584
rect 84244 450400 84564 450720
rect 510000 450240 510320 450560
rect 515564 447560 515884 447880
rect 510660 447240 510980 447560
rect 139640 408673 140640 409673
rect 454544 407060 455544 408060
rect 141040 405673 142040 406673
rect 453144 188447 454144 189447
rect 139640 187060 140640 188060
rect 454544 185447 455544 186447
rect 84244 147560 84564 147880
rect 79236 147240 79556 147560
rect 84904 144560 85224 144880
rect 510660 144400 510980 144720
rect 188447 141488 189447 142488
rect 185447 140088 186447 141088
rect 123400 138556 123720 138876
rect 76236 127240 76556 127560
rect 144400 84244 144720 84564
rect 407060 140088 408060 141088
rect 456460 123400 456780 123720
rect 450240 85690 450560 86010
rect 447240 85030 447560 85350
rect 447560 79236 447880 79556
rect 467560 76236 467880 76556
<< metal3 >>
rect 127240 518884 127560 518894
rect 120560 518564 127240 518884
rect 120560 455448 120880 518564
rect 127240 518554 127560 518564
rect 147240 515884 147560 515894
rect 123560 515564 147240 515884
rect 123560 456108 123880 515564
rect 147240 515554 147560 515564
rect 147560 510532 147880 510541
rect 450400 510532 450720 510541
rect 147551 510212 147560 510532
rect 147880 510212 147889 510532
rect 450391 510212 450400 510532
rect 450720 510212 450729 510532
rect 147560 510203 147880 510212
rect 450400 510203 450720 510212
rect 144560 509872 144880 509881
rect 144551 509552 144560 509872
rect 144880 509552 144889 509872
rect 144560 509543 144880 509552
rect 455800 474560 456120 474570
rect 456120 474240 518884 474560
rect 455800 474230 456120 474240
rect 138444 471720 138764 471729
rect 138435 471400 138444 471720
rect 138764 471400 138773 471720
rect 456460 471560 456780 471570
rect 138444 471391 138764 471400
rect 456780 471240 515884 471560
rect 456460 471230 456780 471240
rect 471400 456332 471720 456341
rect 123550 455788 123560 456108
rect 123880 455788 123890 456108
rect 471391 456012 471400 456332
rect 471720 456012 471729 456332
rect 471400 456003 471720 456012
rect 120550 455128 120560 455448
rect 120880 455128 120890 455448
rect 187060 454984 188060 454993
rect 408673 454984 409673 454993
rect 187051 453984 187060 454984
rect 188060 453984 188069 454984
rect 408664 453984 408673 454984
rect 409673 453984 409682 454984
rect 187060 453975 188060 453984
rect 408673 453975 409673 453984
rect 405673 453584 406673 453593
rect 405664 452584 405673 453584
rect 406673 452584 406682 453584
rect 405673 452575 406673 452584
rect 84244 450720 84564 450729
rect 84235 450400 84244 450720
rect 84564 450400 84573 450720
rect 510000 450560 510320 450569
rect 84244 450391 84564 450400
rect 509991 450240 510000 450560
rect 510320 450240 510329 450560
rect 510000 450231 510320 450240
rect 515564 447880 515884 471240
rect 518564 467880 518884 474240
rect 518554 467560 518564 467880
rect 518884 467560 518894 467880
rect 510660 447560 510980 447569
rect 515554 447560 515564 447880
rect 515884 447560 515894 447880
rect 510651 447240 510660 447560
rect 510980 447240 510989 447560
rect 510660 447231 510980 447240
rect 139640 409673 140640 409682
rect 139631 408673 139640 409673
rect 140640 408673 140649 409673
rect 139640 408664 140640 408673
rect 454544 408060 455544 408069
rect 454535 407060 454544 408060
rect 455544 407060 455553 408060
rect 454544 407051 455544 407060
rect 141040 406673 142040 406682
rect 141031 405673 141040 406673
rect 142040 405673 142049 406673
rect 141040 405664 142040 405673
rect 453144 189447 454144 189456
rect 453135 188447 453144 189447
rect 454144 188447 454153 189447
rect 453144 188438 454144 188447
rect 139640 188060 140640 188069
rect 139631 187060 139640 188060
rect 140640 187060 140649 188060
rect 139640 187051 140640 187060
rect 454544 186447 455544 186456
rect 454535 185447 454544 186447
rect 455544 185447 455553 186447
rect 454544 185438 455544 185447
rect 84244 147880 84564 147889
rect 84235 147560 84244 147880
rect 84564 147560 84573 147880
rect 79226 147240 79236 147560
rect 79556 147240 79566 147560
rect 84244 147551 84564 147560
rect 76226 127240 76236 127560
rect 76556 127240 76566 127560
rect 76236 120880 76556 127240
rect 79236 123880 79556 147240
rect 84904 144880 85224 144889
rect 84895 144560 84904 144880
rect 85224 144560 85233 144880
rect 510660 144720 510980 144729
rect 84904 144551 85224 144560
rect 510651 144400 510660 144720
rect 510980 144400 510989 144720
rect 510660 144391 510980 144400
rect 188447 142488 189447 142497
rect 188438 141488 188447 142488
rect 189447 141488 189456 142488
rect 188447 141479 189447 141488
rect 185447 141088 186447 141097
rect 407060 141088 408060 141097
rect 185438 140088 185447 141088
rect 186447 140088 186456 141088
rect 407051 140088 407060 141088
rect 408060 140088 408069 141088
rect 185447 140079 186447 140088
rect 407060 140079 408060 140088
rect 474230 139400 474240 139720
rect 474560 139400 474570 139720
rect 123400 138876 123720 138885
rect 123391 138556 123400 138876
rect 123720 138556 123729 138876
rect 471230 138740 471240 139060
rect 471560 138740 471570 139060
rect 123400 138547 123720 138556
rect 138444 123880 138764 123890
rect 79236 123560 138444 123880
rect 456460 123720 456780 123729
rect 138444 123550 138764 123560
rect 456451 123400 456460 123720
rect 456780 123400 456789 123720
rect 456460 123391 456780 123400
rect 139104 120880 139424 120890
rect 76236 120560 139104 120880
rect 139104 120550 139424 120560
rect 450240 86010 450560 86019
rect 450231 85690 450240 86010
rect 450560 85690 450569 86010
rect 450240 85681 450560 85690
rect 447240 85350 447560 85359
rect 447231 85030 447240 85350
rect 447560 85030 447569 85350
rect 447240 85021 447560 85030
rect 144400 84564 144720 84573
rect 144391 84244 144400 84564
rect 144720 84244 144729 84564
rect 144400 84235 144720 84244
rect 447560 79556 447880 79566
rect 471240 79556 471560 138740
rect 447880 79236 471560 79556
rect 447560 79226 447880 79236
rect 467560 76556 467880 76566
rect 474240 76556 474560 139400
rect 467880 76236 474560 76556
rect 467560 76226 467880 76236
<< via3 >>
rect 147560 510212 147880 510532
rect 450400 510212 450720 510532
rect 144560 509552 144880 509872
rect 455800 474240 456120 474560
rect 138444 471400 138764 471720
rect 456460 471240 456780 471560
rect 123560 455788 123880 456108
rect 471400 456012 471720 456332
rect 120560 455128 120880 455448
rect 187060 453984 188060 454984
rect 408673 453984 409673 454984
rect 405673 452584 406673 453584
rect 84244 450400 84564 450720
rect 510000 450240 510320 450560
rect 510660 447240 510980 447560
rect 139640 408673 140640 409673
rect 454544 407060 455544 408060
rect 141040 405673 142040 406673
rect 453144 188447 454144 189447
rect 139640 187060 140640 188060
rect 454544 185447 455544 186447
rect 84244 147560 84564 147880
rect 84904 144560 85224 144880
rect 510660 144400 510980 144720
rect 188447 141488 189447 142488
rect 185447 140088 186447 141088
rect 407060 140088 408060 141088
rect 474240 139400 474560 139720
rect 123400 138556 123720 138876
rect 471240 138740 471560 139060
rect 138444 123560 138764 123880
rect 456460 123400 456780 123720
rect 139104 120560 139424 120880
rect 450240 85690 450560 86010
rect 447240 85030 447560 85350
rect 144400 84244 144720 84564
<< metal4 >>
rect 147560 510532 147880 510541
rect 450400 510532 450720 510541
rect 147551 510212 147560 510532
rect 147880 510212 147889 510532
rect 450391 510212 450400 510532
rect 450720 510212 450729 510532
rect 147560 510203 147880 510212
rect 450400 510203 450720 510212
rect 144560 509872 144880 509881
rect 144551 509552 144560 509872
rect 144880 509552 144889 509872
rect 144560 509543 144880 509552
rect 455800 474560 456120 475840
rect 455791 474240 455800 474560
rect 456120 474240 456129 474560
rect 138444 471720 138764 473000
rect 138435 471400 138444 471720
rect 138764 471400 138773 471720
rect 138444 470120 138764 471400
rect 455800 469960 456120 474240
rect 456460 471560 456780 475840
rect 456451 471240 456460 471560
rect 456780 471240 456789 471560
rect 456460 469960 456780 471240
rect 471400 456332 471720 456341
rect 123560 456108 123880 456117
rect 123551 455788 123560 456108
rect 123880 455788 123889 456108
rect 471391 456012 471400 456332
rect 471720 456012 471729 456332
rect 471400 456003 471720 456012
rect 123560 455779 123880 455788
rect 120560 455448 120880 455457
rect 120551 455128 120560 455448
rect 120880 455128 120889 455448
rect 120560 455119 120880 455128
rect 187060 454984 188060 454993
rect 408673 454984 409673 454993
rect 187051 453984 187060 454984
rect 188060 453984 188069 454984
rect 408664 453984 408673 454984
rect 409673 453984 409682 454984
rect 187060 453975 188060 453984
rect 408673 453975 409673 453984
rect 405673 453584 406673 453593
rect 405664 452584 405673 453584
rect 406673 452584 406682 453584
rect 405673 452575 406673 452584
rect 84244 450720 84564 452000
rect 84235 450400 84244 450720
rect 84564 450400 84573 450720
rect 510000 450560 510320 451840
rect 84244 449120 84564 450400
rect 509991 450240 510000 450560
rect 510320 450240 510329 450560
rect 510000 445960 510320 450240
rect 510660 447560 510980 451840
rect 510651 447240 510660 447560
rect 510980 447240 510989 447560
rect 510660 445960 510980 447240
rect 139640 409673 140640 413673
rect 139631 408673 139640 409673
rect 140640 408673 140649 409673
rect 139640 401673 140640 408673
rect 141040 406673 142040 413673
rect 454544 408060 455544 412060
rect 454535 407060 454544 408060
rect 455544 407060 455553 408060
rect 141031 405673 141040 406673
rect 142040 405673 142049 406673
rect 141040 401673 142040 405673
rect 454544 403060 455544 407060
rect 139640 188060 140640 192060
rect 453144 189447 454144 193447
rect 453135 188447 453144 189447
rect 454144 188447 454153 189447
rect 139631 187060 139640 188060
rect 140640 187060 140649 188060
rect 139640 183060 140640 187060
rect 453144 181447 454144 188447
rect 454544 186447 455544 193447
rect 454535 185447 454544 186447
rect 455544 185447 455553 186447
rect 454544 181447 455544 185447
rect 84244 147880 84564 149160
rect 84235 147560 84244 147880
rect 84564 147560 84573 147880
rect 84244 143280 84564 147560
rect 84904 144880 85224 149160
rect 84895 144560 84904 144880
rect 85224 144560 85233 144880
rect 510660 144720 510980 146000
rect 84904 143280 85224 144560
rect 510651 144400 510660 144720
rect 510980 144400 510989 144720
rect 510660 143120 510980 144400
rect 188447 142488 189447 142497
rect 188438 141488 188447 142488
rect 189447 141488 189456 142488
rect 188447 141479 189447 141488
rect 185447 141088 186447 141097
rect 407060 141088 408060 141097
rect 185438 140088 185447 141088
rect 186447 140088 186456 141088
rect 407051 140088 407060 141088
rect 408060 140088 408069 141088
rect 185447 140079 186447 140088
rect 407060 140079 408060 140088
rect 474240 139720 474560 139729
rect 474231 139400 474240 139720
rect 474560 139400 474569 139720
rect 474240 139391 474560 139400
rect 471240 139060 471560 139069
rect 123400 138876 123720 138885
rect 123391 138556 123400 138876
rect 123720 138556 123729 138876
rect 471231 138740 471240 139060
rect 471560 138740 471569 139060
rect 471240 138731 471560 138740
rect 123400 138547 123720 138556
rect 138444 123880 138764 125160
rect 138435 123560 138444 123880
rect 138764 123560 138773 123880
rect 138444 119280 138764 123560
rect 139104 120880 139424 125160
rect 456460 123720 456780 125000
rect 456451 123400 456460 123720
rect 456780 123400 456789 123720
rect 456460 122120 456780 123400
rect 139095 120560 139104 120880
rect 139424 120560 139433 120880
rect 139104 119280 139424 120560
rect 450240 86010 450560 86019
rect 450231 85690 450240 86010
rect 450560 85690 450569 86010
rect 450240 85681 450560 85690
rect 447240 85350 447560 85359
rect 447231 85030 447240 85350
rect 447560 85030 447569 85350
rect 447240 85021 447560 85030
rect 144400 84564 144720 84573
rect 144391 84244 144400 84564
rect 144720 84244 144729 84564
rect 144400 84235 144720 84244
<< via4 >>
rect 147560 510212 147880 510532
rect 450400 510212 450720 510532
rect 144560 509552 144880 509872
rect 123560 455788 123880 456108
rect 471400 456012 471720 456332
rect 120560 455128 120880 455448
rect 187060 453984 188060 454984
rect 408673 453984 409673 454984
rect 405673 452584 406673 453584
rect 188447 141488 189447 142488
rect 185447 140088 186447 141088
rect 407060 140088 408060 141088
rect 474240 139400 474560 139720
rect 123400 138556 123720 138876
rect 471240 138740 471560 139060
rect 450240 85690 450560 86010
rect 447240 85030 447560 85350
rect 144400 84244 144720 84564
<< metal5 >>
rect 147560 510532 147880 510541
rect 450400 510532 450720 510541
rect 143280 510212 147560 510532
rect 147880 510212 149160 510532
rect 449120 510212 450400 510532
rect 450720 510212 452000 510532
rect 147560 510203 147880 510212
rect 450400 510203 450720 510212
rect 144560 509872 144880 509881
rect 143280 509552 144560 509872
rect 144880 509552 149160 509872
rect 144560 509543 144880 509552
rect 471400 456332 471720 456341
rect 123560 456108 123880 456117
rect 119280 455788 123560 456108
rect 123880 455788 125160 456108
rect 470120 456012 471400 456332
rect 471720 456012 473000 456332
rect 471400 456003 471720 456012
rect 123560 455779 123880 455788
rect 120560 455448 120880 455457
rect 119280 455128 120560 455448
rect 120880 455128 125160 455448
rect 120560 455119 120880 455128
rect 187060 454984 188060 454993
rect 408673 454984 409673 454993
rect 183060 453984 187060 454984
rect 188060 453984 192060 454984
rect 401673 453984 408673 454984
rect 409673 453984 413673 454984
rect 187060 453975 188060 453984
rect 408673 453975 409673 453984
rect 405673 453584 406673 453593
rect 401673 452584 405673 453584
rect 406673 452584 413673 453584
rect 405673 452575 406673 452584
rect 188447 142488 189447 142497
rect 181447 141488 188447 142488
rect 189447 141488 193447 142488
rect 188447 141479 189447 141488
rect 185447 141088 186447 141097
rect 407060 141088 408060 141097
rect 181447 140088 185447 141088
rect 186447 140088 193447 141088
rect 403060 140088 407060 141088
rect 408060 140088 412060 141088
rect 185447 140079 186447 140088
rect 407060 140079 408060 140088
rect 474240 139720 474560 139729
rect 469960 139400 474240 139720
rect 474560 139400 475840 139720
rect 474240 139391 474560 139400
rect 471240 139060 471560 139069
rect 123400 138876 123720 138885
rect 122120 138556 123400 138876
rect 123720 138556 125000 138876
rect 469960 138740 471240 139060
rect 471560 138740 475840 139060
rect 471240 138731 471560 138740
rect 123400 138547 123720 138556
rect 450240 86010 450560 86019
rect 445960 85690 450240 86010
rect 450560 85690 451840 86010
rect 450240 85681 450560 85690
rect 447240 85350 447560 85359
rect 445960 85030 447240 85350
rect 447560 85030 451840 85350
rect 447240 85021 447560 85030
rect 144400 84564 144720 84573
rect 143120 84244 144400 84564
rect 144720 84244 146000 84564
rect 144400 84235 144720 84244
use power_taper  power_taper_0
timestamp 1757356513
transform 1 0 120332 0 1 74060
box 0 -200 14456 1344
use power_taper  power_taper_2
timestamp 1757356513
transform 1 0 160332 0 1 74060
box 0 -200 14456 1344
use power_taper  power_taper_3
timestamp 1757356513
transform 1 0 180332 0 1 74060
box 0 -200 14456 1344
use power_taper  power_taper_4
timestamp 1757356513
transform 1 0 400332 0 1 74060
box 0 -200 14456 1344
use power_taper  power_taper_6
timestamp 1757356513
transform 1 0 440332 0 1 74060
box 0 -200 14456 1344
use power_taper  power_taper_7
timestamp 1757356513
transform 1 0 460332 0 1 74060
box 0 -200 14456 1344
use power_taper  power_taper_8
timestamp 1757356513
transform 0 -1 521060 1 0 120332
box 0 -200 14456 1344
use power_taper  power_taper_10
timestamp 1757356513
transform 0 -1 521060 1 0 160332
box 0 -200 14456 1344
use power_taper  power_taper_11
timestamp 1757356513
transform 0 -1 521060 1 0 180332
box 0 -200 14456 1344
use power_taper  power_taper_12
timestamp 1757356513
transform 0 -1 521060 1 0 400332
box 0 -200 14456 1344
use power_taper  power_taper_14
timestamp 1757356513
transform 0 -1 521060 1 0 440332
box 0 -200 14456 1344
use power_taper  power_taper_15
timestamp 1757356513
transform 0 -1 521060 1 0 460332
box 0 -200 14456 1344
use power_taper  power_taper_16
timestamp 1757356513
transform -1 0 474788 0 -1 521060
box 0 -200 14456 1344
use power_taper  power_taper_18
timestamp 1757356513
transform -1 0 434788 0 -1 521060
box 0 -200 14456 1344
use power_taper  power_taper_19
timestamp 1757356513
transform -1 0 414788 0 -1 521060
box 0 -200 14456 1344
use power_taper  power_taper_20
timestamp 1757356513
transform -1 0 194788 0 -1 521060
box 0 -200 14456 1344
use power_taper  power_taper_22
timestamp 1757356513
transform -1 0 154788 0 -1 521060
box 0 -200 14456 1344
use power_taper  power_taper_23
timestamp 1757356513
transform -1 0 134788 0 -1 521060
box 0 -200 14456 1344
use power_taper  power_taper_24
timestamp 1757356513
transform 0 1 74060 -1 0 474788
box 0 -200 14456 1344
use power_taper  power_taper_26
timestamp 1757356513
transform 0 1 74060 -1 0 434788
box 0 -200 14456 1344
use power_taper  power_taper_27
timestamp 1757356513
transform 0 1 74060 -1 0 414788
box 0 -200 14456 1344
use power_taper  power_taper_28
timestamp 1757356513
transform 0 1 74060 -1 0 194788
box 0 -200 14456 1344
use power_taper  power_taper_30
timestamp 1757356513
transform 0 1 74060 -1 0 154788
box 0 -200 14456 1344
use power_taper  power_taper_31
timestamp 1757356513
transform 0 1 74060 -1 0 134788
box 0 -200 14456 1344
use signal_taper  signal_taper_0
timestamp 1757356446
transform 1 0 203128 0 1 74060
box 0 -200 8864 1232
use signal_taper  signal_taper_1
timestamp 1757356446
transform 1 0 223128 0 1 74060
box 0 -200 8864 1232
use signal_taper  signal_taper_2
timestamp 1757356446
transform -1 0 271992 0 -1 521060
box 0 -200 8864 1232
use signal_taper  signal_taper_3
timestamp 1757356446
transform -1 0 251992 0 -1 521060
box 0 -200 8864 1232
use signal_taper  signal_taper_4
timestamp 1757356446
transform -1 0 231992 0 -1 521060
box 0 -200 8864 1232
use signal_taper  signal_taper_5
timestamp 1757356446
transform -1 0 211992 0 -1 521060
box 0 -200 8864 1232
<< labels >>
flabel metal5 143120 84244 146000 84564 0 FreeSans 1024 0 0 0 vss_pad_s_2
port 1 nsew ground bidirectional
flabel metal5 181447 140088 193447 141088 0 FreeSans 1024 0 0 0 vss_pad_s_4
port 2 nsew ground bidirectional
flabel metal5 181447 141488 193447 142488 0 FreeSans 1024 0 0 0 vddcore0_pad_s_5
port 3 nsew power bidirectional
flabel metal5 403060 140088 412060 141088 0 FreeSans 1024 0 0 0 vss_pad_s_16
port 4 nsew ground bidirectional
flabel metal4 510660 143120 510980 146000 0 FreeSans 1024 90 0 0 vss_pad_e_2
port 7 nsew ground bidirectional
flabel metal4 454544 181447 455544 193447 0 FreeSans 1024 90 0 0 vss_pad_e_4
port 8 nsew ground bidirectional
flabel metal4 453144 181447 454144 193447 0 FreeSans 1024 90 0 0 vddcore0_pad_e_5
port 9 nsew power bidirectional
flabel metal4 454544 403060 455544 412060 0 FreeSans 1024 90 0 0 vss_pad_e_16
port 10 nsew ground bidirectional
flabel metal5 449120 510212 452000 510532 0 FreeSans 1024 0 0 0 vss_pad_n_2
port 13 nsew ground bidirectional
flabel metal5 401673 453984 413673 454984 0 FreeSans 1024 0 0 0 vss_pad_n_4
port 14 nsew ground bidirectional
flabel metal5 401673 452584 413673 453584 0 FreeSans 1024 0 0 0 vddcore0_pad_n_5
port 15 nsew power bidirectional
flabel metal5 183060 453984 192060 454984 0 FreeSans 1024 0 0 0 vss_pad_n_16
port 16 nsew ground bidirectional
flabel metal4 84244 449120 84564 452000 0 FreeSans 1024 90 0 0 vss_pad_w_2
port 19 nsew ground bidirectional
flabel metal4 139640 401673 140640 413673 0 FreeSans 1024 90 0 0 vss_pad_w_4
port 20 nsew ground bidirectional
flabel metal4 141040 401673 142040 413673 0 FreeSans 1024 90 0 0 vddcore0_pad_w_5
port 21 nsew power bidirectional
flabel metal4 139640 183060 140640 192060 0 FreeSans 1024 90 0 0 vss_pad_w_16
port 22 nsew ground bidirectional
flabel metal2 207522 75180 207598 76136 0 FreeSans 1024 0 0 0 loop_pad_s_6
port 25 nsew signal bidirectional
flabel metal2 227522 75180 227598 76136 0 FreeSans 1024 0 0 0 loop_pad_s_7
port 26 nsew signal bidirectional
flabel metal2 267522 519384 267598 519940 0 FreeSans 1024 0 0 0 tie_pad_n_12
port 27 nsew signal bidirectional
flabel metal2 247522 518984 247598 519940 0 FreeSans 1024 0 0 0 ta_pad_n_13
port 28 nsew signal bidirectional
flabel metal2 227522 518584 227598 519940 0 FreeSans 1024 0 0 0 toe_pad_n_14
port 29 nsew signal bidirectional
flabel metal2 207522 518184 207598 519940 0 FreeSans 1024 0 0 0 ty_pad_n_15
port 30 nsew signal bidirectional
flabel metal4 84244 143280 84564 149160 0 FreeSans 1024 90 0 0 vss_pad_w_18
port 23 nsew ground bidirectional
flabel metal4 84904 143280 85224 149160 0 FreeSans 1024 90 0 0 vddcore2_pad_w_19
port 24 nsew power bidirectional
flabel metal5 445960 85030 451840 85350 0 FreeSans 1024 0 0 0 vss_pad_s_18
port 5 nsew ground bidirectional
flabel metal5 445960 85690 451840 86010 0 FreeSans 1024 0 0 0 vddcore3_pad_s_19
port 6 nsew power bidirectional
flabel metal4 510660 445960 510980 451840 0 FreeSans 1024 90 0 0 vss_pad_e_18
port 11 nsew ground bidirectional
flabel metal4 510000 445960 510320 451840 0 FreeSans 1024 90 0 0 vddcore4_pad_e_19
port 12 nsew power bidirectional
flabel metal5 143280 510212 149160 510532 0 FreeSans 1024 0 0 0 vss_pad_n_18
port 17 nsew ground bidirectional
flabel metal5 143280 509552 149160 509872 0 FreeSans 1024 0 0 0 vddcore1_pad_n_19
port 18 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 595120 595120
string LEFclass COVER
<< end >>
