magic
tech gf180mcuD
magscale 1 5
timestamp 1757618801
<< metal2 >>
rect 0 0 4432 800
<< end >>
