`default_nettype none

(* blackbox *)
module wiring (
    inout wire vss_pad_s_2,
    inout wire vss_pad_s_4,
    inout wire vddcore0_pad_s_5,
    inout wire vss_pad_s_16,
    inout wire vss_pad_s_18,
    inout wire vddcore3_pad_s_19,
    inout wire vss_pad_e_2,
    inout wire vss_pad_e_4,
    inout wire vddcore0_pad_e_5,
    inout wire vss_pad_e_16,
    inout wire vss_pad_e_18,
    inout wire vddcore4_pad_e_19,
    inout wire vss_pad_n_2,
    inout wire vss_pad_n_4,
    inout wire vddcore0_pad_n_5,
    inout wire vss_pad_n_16,
    inout wire vss_pad_n_18,
    inout wire vddcore1_pad_n_19,
    inout wire vss_pad_w_2,
    inout wire vss_pad_w_4,
    inout wire vddcore0_pad_w_5,
    inout wire vss_pad_w_16,
    inout wire vss_pad_w_18,
    inout wire vddcore2_pad_w_19,
    inout wire loop_pad_s_6,
    inout wire loop_pad_s_7
);

endmodule
