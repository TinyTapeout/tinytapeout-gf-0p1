VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO loopback
  CLASS COVER ;
  FOREIGN loopback ;
  ORIGIN 0.000 0.000 ;
  SIZE 125.000 BY 35.000 ;
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 0.000 25.000 35.000 ;
    END
  END A
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 100.000 0.000 125.000 35.000 ;
    END
  END B
  OBS
      LAYER Metal2 ;
        RECT 25.000 10.000 100.000 35.000 ;
  END
END loopback
END LIBRARY

