magic
tech gf180mcuD
timestamp 1758675408
<< metal2 >>
rect 0 200 2500 700
rect 0 0 500 200
rect 2000 0 2500 200
<< labels >>
flabel metal2 0 0 500 700 0 FreeSans 204 0 0 0 A
port 1 nsew signal bidirectional
flabel metal2 2000 0 2500 700 0 FreeSans 204 0 0 0 B
port 2 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 2500 700
string LEFclass COVER
<< end >>
