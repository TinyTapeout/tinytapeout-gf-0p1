magic
tech gf180mcuD
magscale 1 5
timestamp 1757356513
<< metal2 >>
rect 3600 644 3628 672
rect 3599 616 3629 644
rect 3594 588 3634 616
rect 3589 560 3639 588
rect 3582 532 3646 560
rect 3573 504 3655 532
rect 3561 476 3667 504
rect 3546 448 3682 476
rect 3527 420 3701 448
rect 3503 392 3725 420
rect 3469 364 3759 392
rect 3431 336 3797 364
rect 3379 308 3849 336
rect 3313 280 3915 308
rect 3228 252 4000 280
rect 3119 224 4109 252
rect 2979 196 4249 224
rect 2800 168 4428 196
rect 2571 140 4657 168
rect 2276 112 4952 140
rect 1899 84 5329 112
rect 1415 56 5813 84
rect 795 28 6433 56
rect 0 0 7228 28
use power_conn  power_conn_0
timestamp 1757356272
transform 1 0 -136 0 1 -35000
box 136 34900 7364 35000
<< end >>
