magic
tech gf180mcuD
magscale 1 5
timestamp 1757368090
<< metal2 >>
rect 0 0 14432 4432
<< labels >>
flabel metal2 0 0 4432 4432 0 FreeSans 1024 0 0 0 A
port 1 nsew signal bidirectional
flabel metal2 10000 0 14432 4432 0 FreeSans 1024 0 0 0 B
port 2 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 14432 4432
string LEFclass COVER
<< end >>
