magic
tech gf180mcuD
magscale 1 5
timestamp 1757618869
use power_pad_pin  power_pad_pin_0
timestamp 1757356272
transform 1 0 -136 0 1 -35000
box 136 34900 7364 35000
use power_stub  power_stub_0
timestamp 1757618779
transform 1 0 0 0 1 0
box 0 0 7228 800
use power_taper  power_taper_0
timestamp 1757356513
transform 1 0 0 0 1 800
box 0 0 7228 672
<< end >>
