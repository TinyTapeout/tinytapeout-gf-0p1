magic
tech gf180mcuD
magscale 1 5
timestamp 1757368090
<< metal2 >>
rect 0 0 10038 38
<< labels >>
flabel metal2 0 0 38 38 0 FreeSans 128 0 0 0 A
port 1 nsew signal bidirectional
flabel metal2 10000 0 10038 38 0 FreeSans 128 0 0 0 B
port 2 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 10038 38
string LEFclass COVER
<< end >>
