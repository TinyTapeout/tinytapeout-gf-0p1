VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_logo
  CLASS COVER ;
  FOREIGN tt_logo ;
  ORIGIN 0.000 0.000 ;
  SIZE 225.000 BY 225.000 ;
  PIN dummy
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 105.120 212.040 120.240 212.400 ;
        RECT 101.160 211.680 123.840 212.040 ;
        RECT 98.280 211.320 126.720 211.680 ;
        RECT 95.760 210.960 129.240 211.320 ;
        RECT 93.960 210.600 131.040 210.960 ;
        RECT 92.160 210.240 132.840 210.600 ;
        RECT 90.360 209.880 134.640 210.240 ;
        RECT 88.920 209.520 136.080 209.880 ;
        RECT 87.480 209.160 137.520 209.520 ;
        RECT 86.040 208.800 138.960 209.160 ;
        RECT 84.600 208.440 140.400 208.800 ;
        RECT 83.520 208.080 141.480 208.440 ;
        RECT 82.440 207.720 142.560 208.080 ;
        RECT 81.360 207.360 143.640 207.720 ;
        RECT 80.280 207.000 144.720 207.360 ;
        RECT 79.200 206.640 145.800 207.000 ;
        RECT 78.120 206.280 146.880 206.640 ;
        RECT 77.040 205.920 147.960 206.280 ;
        RECT 76.320 205.560 148.680 205.920 ;
        RECT 75.240 205.200 149.760 205.560 ;
        RECT 74.520 204.840 150.480 205.200 ;
        RECT 73.440 204.480 151.560 204.840 ;
        RECT 72.720 204.120 152.280 204.480 ;
        RECT 72.000 203.760 153.000 204.120 ;
        RECT 70.920 203.400 153.720 203.760 ;
        RECT 70.200 203.040 154.800 203.400 ;
        RECT 69.480 202.680 155.520 203.040 ;
        RECT 68.760 202.320 156.240 202.680 ;
        RECT 68.040 201.960 156.960 202.320 ;
        RECT 67.320 201.600 157.680 201.960 ;
        RECT 66.600 201.240 158.400 201.600 ;
        RECT 65.880 200.880 159.120 201.240 ;
        RECT 65.160 200.520 159.840 200.880 ;
        RECT 64.800 200.160 160.200 200.520 ;
        RECT 64.080 199.800 160.920 200.160 ;
        RECT 63.360 199.440 161.640 199.800 ;
        RECT 62.640 199.080 162.360 199.440 ;
        RECT 61.920 198.720 163.080 199.080 ;
        RECT 61.560 198.360 163.440 198.720 ;
        RECT 60.840 198.000 164.160 198.360 ;
        RECT 60.120 197.640 164.880 198.000 ;
        RECT 59.760 197.280 165.240 197.640 ;
        RECT 59.040 196.920 165.960 197.280 ;
        RECT 58.680 196.560 106.920 196.920 ;
        RECT 118.080 196.560 166.320 196.920 ;
        RECT 57.960 196.200 102.960 196.560 ;
        RECT 122.040 196.200 167.040 196.560 ;
        RECT 57.600 195.840 100.440 196.200 ;
        RECT 124.560 195.840 167.400 196.200 ;
        RECT 56.880 195.480 97.920 195.840 ;
        RECT 127.080 195.480 168.120 195.840 ;
        RECT 56.520 195.120 96.120 195.480 ;
        RECT 128.880 195.120 168.480 195.480 ;
        RECT 55.800 194.760 94.320 195.120 ;
        RECT 130.680 194.760 169.200 195.120 ;
        RECT 55.440 194.400 92.880 194.760 ;
        RECT 132.120 194.400 169.560 194.760 ;
        RECT 54.720 194.040 91.440 194.400 ;
        RECT 133.560 194.040 170.280 194.400 ;
        RECT 54.360 193.680 90.000 194.040 ;
        RECT 135.000 193.680 170.640 194.040 ;
        RECT 53.640 193.320 88.920 193.680 ;
        RECT 136.080 193.320 171.360 193.680 ;
        RECT 53.280 192.960 87.480 193.320 ;
        RECT 137.520 192.960 171.720 193.320 ;
        RECT 52.920 192.600 86.400 192.960 ;
        RECT 138.600 192.600 172.080 192.960 ;
        RECT 52.200 192.240 85.320 192.600 ;
        RECT 139.680 192.240 172.800 192.600 ;
        RECT 51.840 191.880 84.240 192.240 ;
        RECT 140.760 191.880 173.160 192.240 ;
        RECT 51.480 191.520 83.520 191.880 ;
        RECT 141.480 191.520 173.520 191.880 ;
        RECT 51.120 191.160 82.440 191.520 ;
        RECT 142.560 191.160 174.240 191.520 ;
        RECT 50.400 190.800 81.720 191.160 ;
        RECT 143.280 190.800 174.600 191.160 ;
        RECT 50.040 190.440 80.640 190.800 ;
        RECT 144.360 190.440 174.960 190.800 ;
        RECT 49.680 190.080 79.920 190.440 ;
        RECT 145.440 190.080 175.320 190.440 ;
        RECT 48.960 189.720 78.840 190.080 ;
        RECT 146.160 189.720 175.680 190.080 ;
        RECT 48.600 189.360 78.120 189.720 ;
        RECT 146.880 189.360 176.400 189.720 ;
        RECT 48.240 189.000 77.400 189.360 ;
        RECT 147.600 189.000 176.760 189.360 ;
        RECT 47.880 188.640 76.680 189.000 ;
        RECT 148.320 188.640 177.120 189.000 ;
        RECT 47.520 188.280 75.960 188.640 ;
        RECT 149.400 188.280 177.480 188.640 ;
        RECT 47.160 187.920 74.880 188.280 ;
        RECT 149.760 187.920 177.840 188.280 ;
        RECT 46.440 187.560 74.520 187.920 ;
        RECT 150.480 187.560 178.560 187.920 ;
        RECT 46.080 187.200 73.800 187.560 ;
        RECT 151.200 187.200 178.920 187.560 ;
        RECT 45.720 186.840 73.080 187.200 ;
        RECT 151.920 186.840 179.280 187.200 ;
        RECT 45.360 186.480 72.360 186.840 ;
        RECT 152.640 186.480 179.640 186.840 ;
        RECT 45.000 186.120 71.640 186.480 ;
        RECT 153.360 186.120 180.000 186.480 ;
        RECT 44.640 185.760 70.920 186.120 ;
        RECT 154.080 185.760 180.360 186.120 ;
        RECT 44.280 185.400 70.560 185.760 ;
        RECT 154.440 185.400 180.720 185.760 ;
        RECT 43.920 185.040 69.840 185.400 ;
        RECT 155.160 185.040 181.080 185.400 ;
        RECT 43.560 184.680 69.120 185.040 ;
        RECT 155.880 184.680 181.440 185.040 ;
        RECT 43.200 184.320 68.760 184.680 ;
        RECT 156.600 184.320 181.800 184.680 ;
        RECT 42.840 183.960 68.040 184.320 ;
        RECT 156.960 183.960 182.160 184.320 ;
        RECT 42.480 183.600 67.320 183.960 ;
        RECT 157.680 183.600 182.520 183.960 ;
        RECT 42.120 183.240 66.960 183.600 ;
        RECT 158.040 183.240 182.880 183.600 ;
        RECT 41.760 182.880 66.240 183.240 ;
        RECT 158.760 182.880 183.240 183.240 ;
        RECT 41.400 182.520 65.880 182.880 ;
        RECT 159.120 182.520 183.600 182.880 ;
        RECT 41.040 182.160 65.160 182.520 ;
        RECT 159.840 182.160 183.960 182.520 ;
        RECT 40.680 181.800 64.800 182.160 ;
        RECT 160.200 181.800 184.320 182.160 ;
        RECT 40.320 181.440 64.080 181.800 ;
        RECT 160.920 181.440 184.680 181.800 ;
        RECT 39.960 181.080 63.720 181.440 ;
        RECT 161.280 181.080 185.040 181.440 ;
        RECT 39.600 180.720 63.360 181.080 ;
        RECT 161.640 180.720 185.400 181.080 ;
        RECT 39.240 180.360 62.640 180.720 ;
        RECT 162.360 180.360 185.760 180.720 ;
        RECT 38.880 180.000 62.280 180.360 ;
        RECT 162.720 180.000 186.120 180.360 ;
        RECT 38.520 179.640 61.560 180.000 ;
        RECT 163.440 179.640 186.480 180.000 ;
        RECT 38.160 179.280 61.200 179.640 ;
        RECT 163.800 179.280 186.840 179.640 ;
        RECT 37.800 178.920 60.840 179.280 ;
        RECT 164.160 178.920 187.200 179.280 ;
        RECT 37.440 178.560 60.480 178.920 ;
        RECT 164.520 178.560 187.560 178.920 ;
        RECT 37.080 178.200 59.760 178.560 ;
        RECT 165.240 178.200 187.920 178.560 ;
        RECT 37.080 177.840 59.400 178.200 ;
        RECT 165.600 177.840 187.920 178.200 ;
        RECT 36.720 177.480 59.040 177.840 ;
        RECT 165.960 177.480 188.280 177.840 ;
        RECT 36.360 177.120 58.680 177.480 ;
        RECT 166.320 177.120 188.640 177.480 ;
        RECT 36.000 176.760 57.960 177.120 ;
        RECT 167.040 176.760 189.000 177.120 ;
        RECT 35.640 176.400 57.600 176.760 ;
        RECT 167.400 176.400 189.360 176.760 ;
        RECT 35.280 176.040 57.240 176.400 ;
        RECT 167.760 176.040 189.720 176.400 ;
        RECT 34.920 175.680 56.880 176.040 ;
        RECT 168.120 175.680 190.080 176.040 ;
        RECT 34.920 175.320 56.520 175.680 ;
        RECT 168.480 175.320 190.080 175.680 ;
        RECT 34.560 174.960 56.160 175.320 ;
        RECT 168.840 174.960 190.440 175.320 ;
        RECT 34.200 174.600 55.800 174.960 ;
        RECT 169.200 174.600 190.800 174.960 ;
        RECT 33.840 174.240 55.440 174.600 ;
        RECT 169.560 174.240 191.160 174.600 ;
        RECT 33.840 173.880 54.720 174.240 ;
        RECT 169.920 173.880 191.520 174.240 ;
        RECT 33.480 173.520 54.360 173.880 ;
        RECT 170.640 173.520 191.520 173.880 ;
        RECT 33.120 173.160 54.000 173.520 ;
        RECT 171.000 173.160 191.880 173.520 ;
        RECT 32.760 172.800 53.640 173.160 ;
        RECT 171.360 172.800 192.240 173.160 ;
        RECT 32.400 172.440 53.280 172.800 ;
        RECT 171.720 172.440 192.600 172.800 ;
        RECT 32.400 172.080 52.920 172.440 ;
        RECT 172.080 172.080 192.600 172.440 ;
        RECT 32.040 171.720 52.560 172.080 ;
        RECT 172.440 171.720 192.960 172.080 ;
        RECT 31.680 171.360 52.200 171.720 ;
        RECT 172.800 171.360 193.320 171.720 ;
        RECT 31.320 171.000 52.200 171.360 ;
        RECT 173.160 171.000 193.680 171.360 ;
        RECT 31.320 170.640 131.400 171.000 ;
        RECT 173.520 170.640 193.680 171.000 ;
        RECT 30.960 170.280 131.400 170.640 ;
        RECT 30.600 169.560 131.400 170.280 ;
        RECT 173.880 170.280 194.040 170.640 ;
        RECT 173.880 169.920 194.400 170.280 ;
        RECT 174.240 169.560 194.400 169.920 ;
        RECT 30.240 169.200 131.400 169.560 ;
        RECT 174.600 169.200 194.760 169.560 ;
        RECT 29.880 168.480 131.400 169.200 ;
        RECT 174.960 168.840 195.120 169.200 ;
        RECT 175.320 168.480 195.120 168.840 ;
        RECT 29.520 168.120 131.400 168.480 ;
        RECT 175.680 168.120 195.480 168.480 ;
        RECT 29.160 167.400 131.400 168.120 ;
        RECT 176.040 167.760 195.840 168.120 ;
        RECT 176.400 167.400 195.840 167.760 ;
        RECT 28.800 167.040 131.400 167.400 ;
        RECT 176.760 167.040 196.200 167.400 ;
        RECT 28.440 166.320 131.400 167.040 ;
        RECT 177.120 166.320 196.560 167.040 ;
        RECT 28.080 165.960 131.400 166.320 ;
        RECT 177.480 165.960 196.920 166.320 ;
        RECT 27.720 165.240 131.400 165.960 ;
        RECT 177.840 165.600 197.280 165.960 ;
        RECT 178.200 165.240 197.280 165.600 ;
        RECT 27.360 164.880 131.400 165.240 ;
        RECT 27.000 164.160 131.400 164.880 ;
        RECT 178.560 164.880 197.640 165.240 ;
        RECT 178.560 164.520 198.000 164.880 ;
        RECT 178.920 164.160 198.000 164.520 ;
        RECT 26.640 163.440 131.400 164.160 ;
        RECT 179.280 163.800 198.360 164.160 ;
        RECT 179.640 163.440 198.360 163.800 ;
        RECT 26.280 163.080 131.400 163.440 ;
        RECT 25.920 162.360 131.400 163.080 ;
        RECT 180.000 163.080 198.720 163.440 ;
        RECT 180.000 162.720 199.080 163.080 ;
        RECT 180.360 162.360 199.080 162.720 ;
        RECT 25.560 161.640 131.400 162.360 ;
        RECT 180.720 161.640 199.440 162.360 ;
        RECT 25.200 160.920 131.400 161.640 ;
        RECT 181.080 161.280 199.800 161.640 ;
        RECT 181.440 160.920 199.800 161.280 ;
        RECT 24.840 160.200 131.400 160.920 ;
        RECT 181.800 160.560 200.160 160.920 ;
        RECT 181.800 160.200 200.520 160.560 ;
        RECT 24.480 159.840 131.400 160.200 ;
        RECT 182.160 159.840 200.520 160.200 ;
        RECT 24.120 159.120 131.400 159.840 ;
        RECT 182.520 159.120 200.880 159.840 ;
        RECT 23.760 158.400 131.400 159.120 ;
        RECT 182.880 158.760 201.240 159.120 ;
        RECT 23.400 157.680 131.400 158.400 ;
        RECT 183.240 158.400 201.240 158.760 ;
        RECT 183.240 158.040 201.600 158.400 ;
        RECT 183.600 157.680 201.600 158.040 ;
        RECT 23.040 156.960 131.400 157.680 ;
        RECT 183.960 156.960 201.960 157.680 ;
        RECT 22.680 156.240 131.400 156.960 ;
        RECT 184.320 156.600 202.320 156.960 ;
        RECT 22.320 155.520 131.400 156.240 ;
        RECT 184.680 156.240 202.320 156.600 ;
        RECT 184.680 155.880 202.680 156.240 ;
        RECT 21.960 154.800 131.400 155.520 ;
        RECT 185.040 155.520 202.680 155.880 ;
        RECT 185.040 155.160 203.040 155.520 ;
        RECT 21.600 154.080 131.400 154.800 ;
        RECT 185.400 154.800 203.040 155.160 ;
        RECT 185.400 154.440 203.400 154.800 ;
        RECT 185.760 154.080 203.400 154.440 ;
        RECT 21.240 153.000 131.400 154.080 ;
        RECT 186.120 153.360 203.760 154.080 ;
        RECT 20.880 152.280 131.400 153.000 ;
        RECT 186.480 153.000 203.760 153.360 ;
        RECT 186.480 152.640 204.120 153.000 ;
        RECT 20.520 151.560 131.400 152.280 ;
        RECT 186.840 152.280 204.120 152.640 ;
        RECT 186.840 151.920 204.480 152.280 ;
        RECT 20.160 150.480 131.400 151.560 ;
        RECT 187.200 151.560 204.480 151.920 ;
        RECT 187.200 151.200 204.840 151.560 ;
        RECT 187.560 150.480 204.840 151.200 ;
        RECT 19.800 149.760 131.400 150.480 ;
        RECT 187.920 149.760 205.200 150.480 ;
        RECT 19.440 148.680 131.400 149.760 ;
        RECT 188.280 149.040 205.560 149.760 ;
        RECT 19.080 147.960 131.400 148.680 ;
        RECT 188.640 148.680 205.560 149.040 ;
        RECT 188.640 148.320 205.920 148.680 ;
        RECT 18.720 146.880 131.400 147.960 ;
        RECT 189.000 147.960 205.920 148.320 ;
        RECT 189.000 147.600 206.280 147.960 ;
        RECT 189.360 146.880 206.280 147.600 ;
        RECT 18.360 145.800 131.400 146.880 ;
        RECT 189.720 146.160 206.640 146.880 ;
        RECT 18.000 144.720 131.400 145.800 ;
        RECT 190.080 145.800 206.640 146.160 ;
        RECT 190.080 145.080 207.000 145.800 ;
        RECT 17.640 143.640 131.400 144.720 ;
        RECT 190.440 144.360 207.360 145.080 ;
        RECT 17.280 143.280 131.400 143.640 ;
        RECT 190.800 144.000 207.360 144.360 ;
        RECT 190.800 143.280 207.720 144.000 ;
        RECT 14.760 133.560 30.960 135.000 ;
        RECT 14.400 132.480 30.600 133.560 ;
        RECT 14.400 131.760 30.240 132.480 ;
        RECT 14.040 130.680 30.240 131.760 ;
        RECT 14.040 129.600 29.880 130.680 ;
        RECT 13.680 129.240 29.880 129.600 ;
        RECT 13.680 127.440 29.520 129.240 ;
        RECT 13.320 127.080 29.520 127.440 ;
        RECT 13.320 124.920 29.160 127.080 ;
        RECT 13.320 124.560 28.800 124.920 ;
        RECT 12.960 122.400 28.800 124.560 ;
        RECT 12.960 121.320 28.440 122.400 ;
        RECT 12.600 118.800 28.440 121.320 ;
        RECT 72.720 121.680 102.600 143.280 ;
        RECT 191.160 142.920 207.720 143.280 ;
        RECT 191.160 142.560 208.080 142.920 ;
        RECT 191.520 141.480 208.080 142.560 ;
        RECT 191.880 140.760 208.440 141.480 ;
        RECT 192.240 140.400 208.440 140.760 ;
        RECT 192.240 139.680 208.800 140.400 ;
        RECT 192.600 138.960 208.800 139.680 ;
        RECT 192.600 138.600 209.160 138.960 ;
        RECT 192.960 137.880 209.160 138.600 ;
        RECT 192.960 137.520 209.520 137.880 ;
        RECT 193.320 136.440 209.520 137.520 ;
        RECT 193.320 136.080 209.880 136.440 ;
        RECT 193.680 135.000 209.880 136.080 ;
        RECT 194.040 133.560 210.240 135.000 ;
        RECT 194.400 133.200 210.240 133.560 ;
        RECT 194.400 132.120 210.600 133.200 ;
        RECT 194.760 131.400 210.600 132.120 ;
        RECT 194.760 130.680 210.960 131.400 ;
        RECT 195.120 129.240 210.960 130.680 ;
        RECT 195.120 128.880 211.320 129.240 ;
        RECT 195.480 127.080 211.320 128.880 ;
        RECT 195.480 126.720 211.680 127.080 ;
        RECT 195.840 124.560 211.680 126.720 ;
        RECT 196.200 122.040 212.040 124.560 ;
        RECT 12.600 105.840 28.080 118.800 ;
        RECT 12.600 104.040 28.440 105.840 ;
        RECT 12.960 102.600 28.440 104.040 ;
        RECT 12.960 100.440 28.800 102.600 ;
        RECT 13.320 99.720 28.800 100.440 ;
        RECT 13.320 97.560 29.160 99.720 ;
        RECT 13.680 95.760 29.520 97.560 ;
        RECT 13.680 95.400 29.880 95.760 ;
        RECT 14.040 94.320 29.880 95.400 ;
        RECT 14.040 93.600 30.240 94.320 ;
        RECT 14.400 92.520 30.240 93.600 ;
        RECT 72.720 93.960 177.840 121.680 ;
        RECT 196.560 120.960 212.040 122.040 ;
        RECT 196.560 117.720 212.400 120.960 ;
        RECT 196.920 106.920 212.400 117.720 ;
        RECT 196.560 104.040 212.400 106.920 ;
        RECT 196.560 102.960 212.040 104.040 ;
        RECT 196.200 100.440 212.040 102.960 ;
        RECT 195.840 97.920 211.680 100.440 ;
        RECT 195.480 97.560 211.680 97.920 ;
        RECT 195.480 96.120 211.320 97.560 ;
        RECT 195.120 95.400 211.320 96.120 ;
        RECT 195.120 94.320 210.960 95.400 ;
        RECT 14.400 91.800 30.600 92.520 ;
        RECT 14.760 91.080 30.600 91.800 ;
        RECT 14.760 90.000 30.960 91.080 ;
        RECT 15.120 88.560 31.320 90.000 ;
        RECT 15.480 87.480 31.680 88.560 ;
        RECT 15.480 87.120 32.040 87.480 ;
        RECT 15.840 86.400 32.040 87.120 ;
        RECT 15.840 85.680 32.400 86.400 ;
        RECT 16.200 85.320 32.400 85.680 ;
        RECT 16.200 84.600 32.760 85.320 ;
        RECT 16.560 84.240 32.760 84.600 ;
        RECT 16.560 83.160 33.120 84.240 ;
        RECT 16.920 82.440 33.480 83.160 ;
        RECT 16.920 82.080 33.840 82.440 ;
        RECT 17.280 81.360 33.840 82.080 ;
        RECT 17.280 81.000 34.200 81.360 ;
        RECT 17.640 80.640 34.200 81.000 ;
        RECT 17.640 79.920 34.560 80.640 ;
        RECT 18.000 79.560 34.560 79.920 ;
        RECT 18.000 78.840 34.920 79.560 ;
        RECT 18.360 78.120 35.280 78.840 ;
        RECT 18.360 77.760 35.640 78.120 ;
        RECT 18.720 77.040 35.640 77.760 ;
        RECT 19.080 76.320 36.000 77.040 ;
        RECT 19.080 75.960 36.360 76.320 ;
        RECT 19.440 75.600 36.360 75.960 ;
        RECT 72.720 75.600 102.600 93.960 ;
        RECT 19.440 75.240 36.720 75.600 ;
        RECT 19.800 74.880 36.720 75.240 ;
        RECT 19.800 74.160 37.080 74.880 ;
        RECT 20.160 73.440 37.440 74.160 ;
        RECT 20.520 72.720 37.800 73.440 ;
        RECT 20.880 72.000 38.160 72.720 ;
        RECT 20.880 71.640 38.520 72.000 ;
        RECT 21.240 70.920 38.880 71.640 ;
        RECT 21.600 70.200 39.240 70.920 ;
        RECT 21.960 69.840 39.600 70.200 ;
        RECT 21.960 69.480 39.960 69.840 ;
        RECT 22.320 69.120 39.960 69.480 ;
        RECT 22.320 68.760 40.320 69.120 ;
        RECT 22.680 68.400 40.320 68.760 ;
        RECT 22.680 68.040 40.680 68.400 ;
        RECT 23.040 67.320 41.040 68.040 ;
        RECT 23.400 66.600 41.400 67.320 ;
        RECT 23.760 66.240 41.760 66.600 ;
        RECT 23.760 65.880 42.120 66.240 ;
        RECT 24.120 65.520 42.120 65.880 ;
        RECT 24.120 65.160 42.480 65.520 ;
        RECT 24.480 64.440 42.840 65.160 ;
        RECT 24.840 64.080 43.200 64.440 ;
        RECT 24.840 63.720 43.560 64.080 ;
        RECT 25.200 63.360 43.920 63.720 ;
        RECT 25.560 63.000 43.920 63.360 ;
        RECT 25.560 62.640 44.280 63.000 ;
        RECT 25.920 61.920 44.640 62.640 ;
        RECT 26.280 61.560 45.000 61.920 ;
        RECT 26.280 61.200 45.360 61.560 ;
        RECT 26.640 60.840 45.720 61.200 ;
        RECT 27.000 60.120 46.080 60.840 ;
        RECT 27.360 59.760 46.440 60.120 ;
        RECT 27.720 59.400 46.800 59.760 ;
        RECT 27.720 59.040 47.160 59.400 ;
        RECT 28.080 58.320 47.520 59.040 ;
        RECT 28.440 57.960 47.880 58.320 ;
        RECT 28.800 57.600 48.240 57.960 ;
        RECT 28.800 57.240 48.600 57.600 ;
        RECT 29.160 56.880 48.960 57.240 ;
        RECT 29.520 56.520 49.320 56.880 ;
        RECT 29.520 56.160 49.680 56.520 ;
        RECT 29.880 55.800 49.680 56.160 ;
        RECT 30.240 55.440 50.040 55.800 ;
        RECT 30.240 55.080 50.400 55.440 ;
        RECT 30.600 54.720 50.760 55.080 ;
        RECT 30.960 54.360 51.120 54.720 ;
        RECT 31.320 54.000 51.480 54.360 ;
        RECT 31.320 53.640 51.840 54.000 ;
        RECT 31.680 53.280 52.200 53.640 ;
        RECT 32.040 52.920 52.560 53.280 ;
        RECT 32.040 52.560 52.920 52.920 ;
        RECT 32.400 52.200 53.280 52.560 ;
        RECT 32.760 51.840 53.640 52.200 ;
        RECT 33.120 51.480 54.000 51.840 ;
        RECT 33.480 51.120 54.360 51.480 ;
        RECT 33.480 50.760 54.720 51.120 ;
        RECT 33.840 50.400 55.080 50.760 ;
        RECT 34.200 50.040 55.440 50.400 ;
        RECT 34.560 49.680 56.160 50.040 ;
        RECT 34.920 49.320 56.520 49.680 ;
        RECT 34.920 48.960 56.880 49.320 ;
        RECT 35.280 48.600 57.240 48.960 ;
        RECT 35.640 48.240 57.600 48.600 ;
        RECT 36.000 47.880 57.960 48.240 ;
        RECT 36.360 47.520 58.320 47.880 ;
        RECT 36.720 47.160 59.040 47.520 ;
        RECT 36.720 46.800 59.400 47.160 ;
        RECT 37.080 46.440 59.760 46.800 ;
        RECT 37.440 46.080 60.120 46.440 ;
        RECT 37.800 45.720 60.840 46.080 ;
        RECT 38.160 45.360 61.200 45.720 ;
        RECT 38.520 45.000 61.560 45.360 ;
        RECT 38.880 44.640 62.280 45.000 ;
        RECT 39.240 44.280 62.640 44.640 ;
        RECT 39.600 43.920 63.000 44.280 ;
        RECT 39.960 43.560 63.720 43.920 ;
        RECT 39.960 43.200 64.080 43.560 ;
        RECT 40.320 42.840 64.800 43.200 ;
        RECT 40.680 42.480 65.160 42.840 ;
        RECT 41.040 42.120 65.520 42.480 ;
        RECT 41.400 41.760 66.240 42.120 ;
        RECT 41.760 41.400 66.960 41.760 ;
        RECT 42.120 41.040 67.320 41.400 ;
        RECT 42.480 40.680 68.040 41.040 ;
        RECT 42.840 40.320 68.400 40.680 ;
        RECT 43.200 39.960 69.120 40.320 ;
        RECT 43.920 39.600 69.840 39.960 ;
        RECT 44.280 39.240 70.200 39.600 ;
        RECT 44.640 38.880 70.920 39.240 ;
        RECT 45.000 38.520 71.640 38.880 ;
        RECT 45.360 38.160 72.360 38.520 ;
        RECT 45.720 37.800 73.080 38.160 ;
        RECT 46.080 37.440 73.800 37.800 ;
        RECT 46.440 37.080 74.160 37.440 ;
        RECT 46.800 36.720 74.880 37.080 ;
        RECT 47.520 36.360 75.600 36.720 ;
        RECT 47.880 36.000 76.320 36.360 ;
        RECT 48.240 35.640 77.400 36.000 ;
        RECT 48.600 35.280 78.120 35.640 ;
        RECT 48.960 34.920 78.840 35.280 ;
        RECT 49.680 34.560 79.560 34.920 ;
        RECT 50.040 34.200 80.640 34.560 ;
        RECT 50.400 33.840 81.360 34.200 ;
        RECT 50.760 33.480 82.440 33.840 ;
        RECT 51.480 33.120 83.160 33.480 ;
        RECT 51.840 32.760 84.240 33.120 ;
        RECT 52.200 32.400 85.320 32.760 ;
        RECT 52.920 32.040 86.400 32.400 ;
        RECT 53.280 31.680 87.480 32.040 ;
        RECT 53.640 31.320 88.920 31.680 ;
        RECT 54.360 30.960 90.000 31.320 ;
        RECT 54.720 30.600 91.440 30.960 ;
        RECT 55.440 30.240 92.880 30.600 ;
        RECT 55.800 29.880 94.320 30.240 ;
        RECT 56.160 29.520 96.120 29.880 ;
        RECT 56.880 29.160 98.280 29.520 ;
        RECT 57.240 28.800 100.080 29.160 ;
        RECT 57.960 28.440 102.960 28.800 ;
        RECT 119.160 28.440 149.040 93.960 ;
        RECT 194.760 93.600 210.960 94.320 ;
        RECT 194.760 92.880 210.600 93.600 ;
        RECT 194.400 91.800 210.600 92.880 ;
        RECT 194.400 91.440 210.240 91.800 ;
        RECT 194.040 90.000 210.240 91.440 ;
        RECT 193.680 88.920 209.880 90.000 ;
        RECT 193.320 88.560 209.880 88.920 ;
        RECT 193.320 87.480 209.520 88.560 ;
        RECT 192.960 87.120 209.520 87.480 ;
        RECT 192.960 86.400 209.160 87.120 ;
        RECT 192.600 85.680 209.160 86.400 ;
        RECT 192.600 85.320 208.800 85.680 ;
        RECT 192.240 84.600 208.800 85.320 ;
        RECT 192.240 84.240 208.440 84.600 ;
        RECT 191.880 83.520 208.440 84.240 ;
        RECT 191.520 83.160 208.440 83.520 ;
        RECT 191.520 82.440 208.080 83.160 ;
        RECT 191.160 82.080 208.080 82.440 ;
        RECT 191.160 81.360 207.720 82.080 ;
        RECT 190.800 81.000 207.720 81.360 ;
        RECT 190.800 80.640 207.360 81.000 ;
        RECT 190.440 79.920 207.360 80.640 ;
        RECT 190.080 78.840 207.000 79.920 ;
        RECT 189.720 78.120 206.640 78.840 ;
        RECT 189.360 77.760 206.640 78.120 ;
        RECT 189.360 77.400 206.280 77.760 ;
        RECT 189.000 77.040 206.280 77.400 ;
        RECT 189.000 76.680 205.920 77.040 ;
        RECT 188.640 75.960 205.920 76.680 ;
        RECT 188.640 75.600 205.560 75.960 ;
        RECT 188.280 75.240 205.560 75.600 ;
        RECT 188.280 74.880 205.200 75.240 ;
        RECT 187.920 74.160 205.200 74.880 ;
        RECT 187.560 73.800 204.840 74.160 ;
        RECT 187.200 73.440 204.840 73.800 ;
        RECT 187.200 73.080 204.480 73.440 ;
        RECT 186.840 72.720 204.480 73.080 ;
        RECT 186.840 72.360 204.120 72.720 ;
        RECT 186.480 71.640 204.120 72.360 ;
        RECT 186.120 70.920 203.760 71.640 ;
        RECT 185.760 70.200 203.400 70.920 ;
        RECT 185.400 69.840 203.040 70.200 ;
        RECT 185.040 69.480 203.040 69.840 ;
        RECT 185.040 69.120 202.680 69.480 ;
        RECT 184.680 68.760 202.680 69.120 ;
        RECT 184.680 68.400 202.320 68.760 ;
        RECT 184.320 68.040 202.320 68.400 ;
        RECT 183.960 67.320 201.960 68.040 ;
        RECT 183.600 66.960 201.600 67.320 ;
        RECT 183.240 66.600 201.600 66.960 ;
        RECT 183.240 66.240 201.240 66.600 ;
        RECT 182.880 65.880 201.240 66.240 ;
        RECT 182.520 65.160 200.880 65.880 ;
        RECT 182.160 64.800 200.520 65.160 ;
        RECT 181.800 64.440 200.520 64.800 ;
        RECT 181.800 64.080 200.160 64.440 ;
        RECT 181.440 63.720 200.160 64.080 ;
        RECT 181.080 63.360 199.800 63.720 ;
        RECT 181.080 63.000 199.440 63.360 ;
        RECT 180.720 62.640 199.440 63.000 ;
        RECT 180.360 62.280 199.080 62.640 ;
        RECT 180.000 61.920 199.080 62.280 ;
        RECT 180.000 61.560 198.720 61.920 ;
        RECT 179.640 61.200 198.720 61.560 ;
        RECT 179.280 60.840 198.360 61.200 ;
        RECT 178.920 60.120 198.000 60.840 ;
        RECT 178.560 59.760 197.640 60.120 ;
        RECT 178.200 59.400 197.640 59.760 ;
        RECT 177.840 59.040 197.280 59.400 ;
        RECT 177.480 58.680 196.920 59.040 ;
        RECT 177.120 58.320 196.920 58.680 ;
        RECT 177.120 57.960 196.560 58.320 ;
        RECT 176.760 57.600 196.200 57.960 ;
        RECT 176.400 57.240 196.200 57.600 ;
        RECT 176.040 56.880 195.840 57.240 ;
        RECT 175.680 56.520 195.480 56.880 ;
        RECT 175.320 56.160 195.480 56.520 ;
        RECT 174.960 55.800 195.120 56.160 ;
        RECT 174.600 55.080 194.760 55.800 ;
        RECT 174.240 54.720 194.400 55.080 ;
        RECT 173.880 54.360 194.040 54.720 ;
        RECT 173.520 54.000 193.680 54.360 ;
        RECT 173.160 53.640 193.680 54.000 ;
        RECT 172.800 53.280 193.320 53.640 ;
        RECT 172.440 52.920 192.960 53.280 ;
        RECT 172.080 52.560 192.960 52.920 ;
        RECT 171.720 52.200 192.600 52.560 ;
        RECT 171.360 51.840 192.240 52.200 ;
        RECT 171.000 51.480 191.880 51.840 ;
        RECT 170.640 51.120 191.880 51.480 ;
        RECT 170.280 50.760 191.520 51.120 ;
        RECT 169.920 50.400 191.160 50.760 ;
        RECT 169.200 50.040 190.800 50.400 ;
        RECT 168.840 49.680 190.440 50.040 ;
        RECT 168.480 49.320 190.440 49.680 ;
        RECT 168.120 48.960 190.080 49.320 ;
        RECT 167.760 48.600 189.720 48.960 ;
        RECT 167.400 48.240 189.360 48.600 ;
        RECT 167.040 47.880 189.000 48.240 ;
        RECT 166.320 47.520 188.640 47.880 ;
        RECT 165.960 47.160 188.640 47.520 ;
        RECT 165.600 46.800 188.280 47.160 ;
        RECT 165.240 46.440 187.920 46.800 ;
        RECT 164.880 46.080 187.560 46.440 ;
        RECT 164.160 45.720 187.200 46.080 ;
        RECT 163.800 45.360 186.840 45.720 ;
        RECT 163.440 45.000 186.480 45.360 ;
        RECT 162.720 44.640 186.120 45.000 ;
        RECT 162.360 44.280 185.760 44.640 ;
        RECT 162.000 43.920 185.400 44.280 ;
        RECT 161.280 43.560 185.400 43.920 ;
        RECT 160.920 43.200 185.040 43.560 ;
        RECT 160.200 42.840 184.680 43.200 ;
        RECT 159.840 42.480 184.320 42.840 ;
        RECT 159.120 42.120 183.960 42.480 ;
        RECT 158.760 41.760 183.600 42.120 ;
        RECT 158.040 41.400 183.240 41.760 ;
        RECT 157.680 41.040 182.880 41.400 ;
        RECT 58.320 28.080 106.920 28.440 ;
        RECT 117.720 28.080 149.040 28.440 ;
        RECT 59.040 27.720 149.040 28.080 ;
        RECT 59.760 27.360 149.040 27.720 ;
        RECT 60.120 27.000 149.040 27.360 ;
        RECT 60.840 26.640 149.040 27.000 ;
        RECT 61.560 26.280 149.040 26.640 ;
        RECT 61.920 25.920 149.040 26.280 ;
        RECT 62.640 25.560 149.040 25.920 ;
        RECT 63.360 25.200 149.040 25.560 ;
        RECT 64.080 24.840 149.040 25.200 ;
        RECT 64.440 24.480 149.040 24.840 ;
        RECT 65.160 24.120 149.040 24.480 ;
        RECT 65.880 23.760 149.040 24.120 ;
        RECT 66.600 23.400 149.040 23.760 ;
        RECT 157.320 40.680 182.520 41.040 ;
        RECT 157.320 40.320 182.160 40.680 ;
        RECT 157.320 39.960 181.800 40.320 ;
        RECT 157.320 39.600 181.440 39.960 ;
        RECT 157.320 39.240 180.720 39.600 ;
        RECT 157.320 38.880 180.360 39.240 ;
        RECT 157.320 38.520 180.000 38.880 ;
        RECT 157.320 38.160 179.640 38.520 ;
        RECT 157.320 37.800 179.280 38.160 ;
        RECT 157.320 37.440 178.920 37.800 ;
        RECT 157.320 37.080 178.560 37.440 ;
        RECT 157.320 36.720 178.200 37.080 ;
        RECT 157.320 36.360 177.840 36.720 ;
        RECT 157.320 36.000 177.120 36.360 ;
        RECT 157.320 35.640 176.760 36.000 ;
        RECT 157.320 35.280 176.400 35.640 ;
        RECT 157.320 34.920 176.040 35.280 ;
        RECT 157.320 34.560 175.680 34.920 ;
        RECT 157.320 34.200 174.960 34.560 ;
        RECT 157.320 33.840 174.600 34.200 ;
        RECT 157.320 33.480 174.240 33.840 ;
        RECT 157.320 33.120 173.520 33.480 ;
        RECT 157.320 32.760 173.160 33.120 ;
        RECT 157.320 32.400 172.800 32.760 ;
        RECT 157.320 32.040 172.440 32.400 ;
        RECT 157.320 31.680 171.720 32.040 ;
        RECT 157.320 31.320 171.360 31.680 ;
        RECT 157.320 30.960 170.640 31.320 ;
        RECT 157.320 30.600 170.280 30.960 ;
        RECT 157.320 30.240 169.920 30.600 ;
        RECT 157.320 29.880 169.200 30.240 ;
        RECT 157.320 29.520 168.840 29.880 ;
        RECT 157.320 29.160 168.120 29.520 ;
        RECT 157.320 28.800 167.760 29.160 ;
        RECT 157.320 28.440 167.040 28.800 ;
        RECT 157.320 28.080 166.680 28.440 ;
        RECT 157.320 27.720 165.960 28.080 ;
        RECT 157.320 27.360 165.600 27.720 ;
        RECT 157.320 27.000 164.880 27.360 ;
        RECT 157.320 26.640 164.160 27.000 ;
        RECT 157.320 26.280 163.800 26.640 ;
        RECT 157.320 25.920 163.080 26.280 ;
        RECT 157.320 25.560 162.360 25.920 ;
        RECT 157.320 25.200 161.640 25.560 ;
        RECT 157.320 24.840 161.280 25.200 ;
        RECT 157.320 24.480 160.560 24.840 ;
        RECT 157.320 24.120 159.840 24.480 ;
        RECT 157.320 23.760 159.120 24.120 ;
        RECT 157.320 23.400 158.400 23.760 ;
        RECT 67.320 23.040 149.040 23.400 ;
        RECT 68.040 22.680 149.040 23.040 ;
        RECT 68.760 22.320 149.040 22.680 ;
        RECT 69.480 21.960 149.040 22.320 ;
        RECT 70.200 21.600 149.040 21.960 ;
        RECT 70.920 21.240 149.040 21.600 ;
        RECT 72.000 20.880 149.040 21.240 ;
        RECT 72.720 20.520 149.040 20.880 ;
        RECT 73.440 20.160 149.040 20.520 ;
        RECT 74.520 19.800 149.040 20.160 ;
        RECT 75.240 19.440 149.040 19.800 ;
        RECT 76.320 19.080 148.680 19.440 ;
        RECT 77.040 18.720 147.960 19.080 ;
        RECT 78.120 18.360 146.880 18.720 ;
        RECT 79.200 18.000 145.800 18.360 ;
        RECT 80.280 17.640 144.720 18.000 ;
        RECT 81.360 17.280 143.640 17.640 ;
        RECT 82.440 16.920 142.560 17.280 ;
        RECT 83.520 16.560 141.480 16.920 ;
        RECT 84.600 16.200 140.400 16.560 ;
        RECT 86.040 15.840 138.960 16.200 ;
        RECT 87.480 15.480 137.520 15.840 ;
        RECT 88.920 15.120 136.080 15.480 ;
        RECT 90.360 14.760 134.640 15.120 ;
        RECT 91.800 14.400 132.840 14.760 ;
        RECT 93.960 14.040 131.040 14.400 ;
        RECT 95.760 13.680 128.880 14.040 ;
        RECT 98.280 13.320 126.720 13.680 ;
        RECT 101.160 12.960 123.840 13.320 ;
        RECT 104.760 12.600 120.240 12.960 ;
    END
  END dummy
END tt_logo
END LIBRARY

